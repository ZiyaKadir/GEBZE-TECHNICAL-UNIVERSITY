magic
tech scmos
timestamp 1736876954
<< nwell >>
rect -78 172 421 200
<< ntransistor >>
rect -67 114 -65 118
rect -59 114 -57 118
rect -43 114 -41 118
rect -27 114 -25 118
rect -10 114 -8 118
rect -4 114 -2 118
rect 28 114 30 118
rect 52 114 54 118
rect 58 114 60 118
rect 76 114 78 118
rect 92 114 94 118
rect 100 114 102 118
rect 116 114 118 118
rect 124 114 126 118
rect 140 114 142 118
rect 148 114 150 118
rect 164 114 166 118
rect 172 114 174 118
rect 189 114 191 118
rect 197 114 199 118
rect 229 114 231 118
rect 235 114 237 118
rect 265 114 267 118
rect 271 114 273 118
rect 289 114 291 118
rect 305 114 307 118
rect 313 114 315 118
rect 329 114 331 118
rect 337 114 339 118
rect 353 114 355 118
rect 361 114 363 118
rect 377 114 379 118
rect 385 114 387 118
rect 402 114 404 118
rect 410 114 412 118
<< ptransistor >>
rect -67 178 -65 186
rect -61 178 -59 186
rect -43 178 -41 186
rect -27 178 -25 186
rect -10 178 -8 186
rect -2 178 0 186
rect 28 178 30 186
rect 52 178 54 186
rect 60 178 62 186
rect 76 178 78 186
rect 92 178 94 186
rect 98 178 100 186
rect 116 178 118 186
rect 122 178 124 186
rect 140 178 142 186
rect 146 178 148 186
rect 164 178 166 186
rect 170 178 172 186
rect 189 178 191 186
rect 195 178 197 186
rect 229 178 231 186
rect 237 178 239 186
rect 265 178 267 186
rect 273 178 275 186
rect 289 178 291 186
rect 305 178 307 186
rect 311 178 313 186
rect 329 178 331 186
rect 335 178 337 186
rect 353 178 355 186
rect 359 178 361 186
rect 377 178 379 186
rect 383 178 385 186
rect 402 178 404 186
rect 408 178 410 186
<< ndiffusion >>
rect -68 114 -67 118
rect -65 114 -64 118
rect -60 114 -59 118
rect -57 114 -56 118
rect -44 114 -43 118
rect -41 114 -40 118
rect -28 114 -27 118
rect -25 114 -24 118
rect -11 114 -10 118
rect -8 114 -4 118
rect -2 114 -1 118
rect 27 114 28 118
rect 30 114 31 118
rect 51 114 52 118
rect 54 114 58 118
rect 60 114 61 118
rect 75 114 76 118
rect 78 114 79 118
rect 91 114 92 118
rect 94 114 95 118
rect 99 114 100 118
rect 102 114 103 118
rect 115 114 116 118
rect 118 114 119 118
rect 123 114 124 118
rect 126 114 127 118
rect 139 114 140 118
rect 142 114 143 118
rect 147 114 148 118
rect 150 114 151 118
rect 163 114 164 118
rect 166 114 167 118
rect 171 114 172 118
rect 174 114 175 118
rect 188 114 189 118
rect 191 114 192 118
rect 196 114 197 118
rect 199 114 200 118
rect 228 114 229 118
rect 231 114 235 118
rect 237 114 238 118
rect 264 114 265 118
rect 267 114 271 118
rect 273 114 274 118
rect 288 114 289 118
rect 291 114 292 118
rect 304 114 305 118
rect 307 114 308 118
rect 312 114 313 118
rect 315 114 316 118
rect 328 114 329 118
rect 331 114 332 118
rect 336 114 337 118
rect 339 114 340 118
rect 352 114 353 118
rect 355 114 356 118
rect 360 114 361 118
rect 363 114 364 118
rect 376 114 377 118
rect 379 114 380 118
rect 384 114 385 118
rect 387 114 388 118
rect 401 114 402 118
rect 404 114 405 118
rect 409 114 410 118
rect 412 114 413 118
<< pdiffusion >>
rect -68 178 -67 186
rect -65 178 -61 186
rect -59 178 -58 186
rect -44 178 -43 186
rect -41 178 -40 186
rect -28 178 -27 186
rect -25 178 -24 186
rect -11 178 -10 186
rect -8 178 -7 186
rect -3 178 -2 186
rect 0 178 1 186
rect 27 178 28 186
rect 30 178 31 186
rect 51 178 52 186
rect 54 178 55 186
rect 59 178 60 186
rect 62 178 63 186
rect 75 178 76 186
rect 78 178 79 186
rect 91 178 92 186
rect 94 178 98 186
rect 100 178 101 186
rect 115 178 116 186
rect 118 178 122 186
rect 124 178 125 186
rect 139 178 140 186
rect 142 178 146 186
rect 148 178 149 186
rect 163 178 164 186
rect 166 178 170 186
rect 172 178 173 186
rect 188 178 189 186
rect 191 178 195 186
rect 197 178 198 186
rect 228 178 229 186
rect 231 178 232 186
rect 236 178 237 186
rect 239 178 240 186
rect 264 178 265 186
rect 267 178 268 186
rect 272 178 273 186
rect 275 178 276 186
rect 288 178 289 186
rect 291 178 292 186
rect 304 178 305 186
rect 307 178 311 186
rect 313 178 314 186
rect 328 178 329 186
rect 331 178 335 186
rect 337 178 338 186
rect 352 178 353 186
rect 355 178 359 186
rect 361 178 362 186
rect 376 178 377 186
rect 379 178 383 186
rect 385 178 386 186
rect 401 178 402 186
rect 404 178 408 186
rect 410 178 411 186
<< ndcontact >>
rect -72 114 -68 118
rect -64 114 -60 118
rect -56 114 -52 118
rect -48 114 -44 118
rect -40 114 -36 118
rect -32 114 -28 118
rect -24 114 -20 118
rect -15 114 -11 118
rect -1 114 3 118
rect 23 114 27 118
rect 31 114 35 118
rect 47 114 51 118
rect 61 114 65 118
rect 71 114 75 118
rect 79 114 83 118
rect 87 114 91 118
rect 95 114 99 118
rect 103 114 107 118
rect 111 114 115 118
rect 119 114 123 118
rect 127 114 131 118
rect 135 114 139 118
rect 143 114 147 118
rect 151 114 155 118
rect 159 114 163 118
rect 167 114 171 118
rect 175 114 179 118
rect 184 114 188 118
rect 192 114 196 118
rect 200 114 204 118
rect 224 114 228 118
rect 238 114 242 118
rect 260 114 264 118
rect 274 114 278 118
rect 284 114 288 118
rect 292 114 296 118
rect 300 114 304 118
rect 308 114 312 118
rect 316 114 320 118
rect 324 114 328 118
rect 332 114 336 118
rect 340 114 344 118
rect 348 114 352 118
rect 356 114 360 118
rect 364 114 368 118
rect 372 114 376 118
rect 380 114 384 118
rect 388 114 392 118
rect 397 114 401 118
rect 405 114 409 118
rect 413 114 417 118
<< pdcontact >>
rect -72 178 -68 186
rect -58 178 -54 186
rect -48 178 -44 186
rect -40 178 -36 186
rect -32 178 -28 186
rect -24 178 -20 186
rect -15 178 -11 186
rect -7 178 -3 186
rect 1 178 5 186
rect 23 178 27 186
rect 31 178 35 186
rect 47 178 51 186
rect 55 178 59 186
rect 63 178 67 186
rect 71 178 75 186
rect 79 178 83 186
rect 87 178 91 186
rect 101 178 105 186
rect 111 178 115 186
rect 125 178 129 186
rect 135 178 139 186
rect 149 178 153 186
rect 159 178 163 186
rect 173 178 177 186
rect 184 178 188 186
rect 198 178 202 186
rect 224 178 228 186
rect 232 178 236 186
rect 240 178 244 186
rect 260 178 264 186
rect 268 178 272 186
rect 276 178 280 186
rect 284 178 288 186
rect 292 178 296 186
rect 300 178 304 186
rect 314 178 318 186
rect 324 178 328 186
rect 338 178 342 186
rect 348 178 352 186
rect 362 178 366 186
rect 372 178 376 186
rect 386 178 390 186
rect 397 178 401 186
rect 411 178 415 186
<< psubstratepcontact >>
rect -72 105 -68 109
rect -64 105 -60 109
rect -56 105 -52 109
rect -48 103 -44 107
rect -40 103 -36 107
rect -32 103 -28 107
rect -24 103 -20 107
rect -15 103 -11 107
rect -4 103 0 107
rect 23 103 27 107
rect 31 103 35 107
rect 47 103 51 107
rect 58 103 62 107
rect 71 103 75 107
rect 79 103 83 107
rect 87 105 91 109
rect 95 105 99 109
rect 103 105 107 109
rect 111 105 115 109
rect 119 105 123 109
rect 127 105 131 109
rect 135 105 139 109
rect 143 105 147 109
rect 151 105 155 109
rect 159 105 163 109
rect 167 105 171 109
rect 175 105 179 109
rect 184 105 188 109
rect 192 105 196 109
rect 200 105 204 109
rect 224 103 228 107
rect 235 103 239 107
rect 260 103 264 107
rect 271 103 275 107
rect 284 103 288 107
rect 292 103 296 107
rect 300 105 304 109
rect 308 105 312 109
rect 316 105 320 109
rect 324 105 328 109
rect 332 105 336 109
rect 340 105 344 109
rect 348 105 352 109
rect 356 105 360 109
rect 364 105 368 109
rect 372 105 376 109
rect 380 105 384 109
rect 388 105 392 109
rect 397 105 401 109
rect 405 105 409 109
rect 413 105 417 109
<< nsubstratencontact >>
rect -72 191 -68 195
rect -58 191 -54 195
rect -48 193 -44 197
rect -40 193 -36 197
rect -32 193 -28 197
rect -24 193 -20 197
rect -15 193 -11 197
rect -7 193 -3 197
rect 1 193 5 197
rect 23 193 27 197
rect 31 193 35 197
rect 47 193 51 197
rect 55 193 59 197
rect 63 193 67 197
rect 71 193 75 197
rect 79 193 83 197
rect 87 191 91 195
rect 101 191 105 195
rect 111 191 115 195
rect 125 191 129 195
rect 135 191 139 195
rect 149 191 153 195
rect 159 191 163 195
rect 173 191 177 195
rect 184 191 188 195
rect 198 191 202 195
rect 224 193 228 197
rect 232 193 236 197
rect 240 193 244 197
rect 260 193 264 197
rect 268 193 272 197
rect 276 193 280 197
rect 284 193 288 197
rect 292 193 296 197
rect 300 191 304 195
rect 314 191 318 195
rect 324 191 328 195
rect 338 191 342 195
rect 348 191 352 195
rect 362 191 366 195
rect 372 191 376 195
rect 386 191 390 195
rect 397 191 401 195
rect 411 191 415 195
<< polysilicon >>
rect -67 186 -65 189
rect -61 186 -59 189
rect -43 186 -41 189
rect -27 186 -25 189
rect -10 186 -8 189
rect -2 186 0 189
rect 28 186 30 189
rect 52 186 54 189
rect 60 186 62 189
rect 76 186 78 189
rect 92 186 94 189
rect 98 186 100 189
rect 116 186 118 189
rect 122 186 124 189
rect 140 186 142 189
rect 146 186 148 189
rect 164 186 166 189
rect 170 186 172 189
rect 189 186 191 189
rect 195 186 197 189
rect 229 186 231 189
rect 237 186 239 189
rect 265 186 267 189
rect 273 186 275 189
rect 289 186 291 189
rect 305 186 307 189
rect 311 186 313 189
rect 329 186 331 189
rect 335 186 337 189
rect 353 186 355 189
rect 359 186 361 189
rect 377 186 379 189
rect 383 186 385 189
rect 402 186 404 189
rect 408 186 410 189
rect -67 118 -65 178
rect -61 177 -59 178
rect -61 175 -57 177
rect -59 118 -57 175
rect -43 118 -41 178
rect -27 118 -25 178
rect -10 118 -8 178
rect -2 122 0 178
rect -4 120 0 122
rect -4 118 -2 120
rect 28 118 30 178
rect 52 118 54 178
rect 60 122 62 178
rect 58 120 62 122
rect 58 118 60 120
rect 76 118 78 178
rect 92 118 94 178
rect 98 177 100 178
rect 98 175 102 177
rect 100 118 102 175
rect 116 118 118 178
rect 122 177 124 178
rect 122 175 126 177
rect 124 118 126 175
rect 140 118 142 178
rect 146 177 148 178
rect 146 175 150 177
rect 148 118 150 175
rect 164 118 166 178
rect 170 177 172 178
rect 170 175 174 177
rect 172 118 174 175
rect 189 118 191 178
rect 195 177 197 178
rect 195 175 199 177
rect 197 118 199 175
rect 229 118 231 178
rect 237 122 239 178
rect 235 120 239 122
rect 235 118 237 120
rect 265 118 267 178
rect 273 122 275 178
rect 271 120 275 122
rect 271 118 273 120
rect 289 118 291 178
rect 305 118 307 178
rect 311 177 313 178
rect 311 175 315 177
rect 313 118 315 175
rect 329 118 331 178
rect 335 177 337 178
rect 335 175 339 177
rect 337 118 339 175
rect 353 118 355 178
rect 359 177 361 178
rect 359 175 363 177
rect 361 118 363 175
rect 377 118 379 178
rect 383 177 385 178
rect 383 175 387 177
rect 385 118 387 175
rect 402 118 404 178
rect 408 177 410 178
rect 408 175 412 177
rect 410 118 412 175
rect -67 111 -65 114
rect -59 111 -57 114
rect -43 111 -41 114
rect -27 111 -25 114
rect -10 111 -8 114
rect -4 111 -2 114
rect 28 111 30 114
rect 52 111 54 114
rect 58 111 60 114
rect 76 111 78 114
rect 92 111 94 114
rect 100 111 102 114
rect 116 111 118 114
rect 124 111 126 114
rect 140 111 142 114
rect 148 111 150 114
rect 164 111 166 114
rect 172 111 174 114
rect 189 111 191 114
rect 197 111 199 114
rect 229 111 231 114
rect 235 111 237 114
rect 265 111 267 114
rect 271 111 273 114
rect 289 111 291 114
rect 305 111 307 114
rect 313 111 315 114
rect 329 111 331 114
rect 337 111 339 114
rect 353 111 355 114
rect 361 111 363 114
rect 377 111 379 114
rect 385 111 387 114
rect 402 111 404 114
rect 410 111 412 114
<< polycontact >>
rect -71 167 -67 171
rect -57 167 -53 171
rect -47 148 -43 152
rect -31 168 -27 172
rect 72 133 76 137
rect 88 121 92 125
rect 136 141 140 145
rect 160 127 164 131
rect 185 166 189 170
rect 285 133 289 137
rect 301 121 305 125
rect 349 121 353 125
rect 373 127 377 131
rect 398 166 402 170
<< metal1 >>
rect -72 197 415 198
rect -72 195 -48 197
rect -68 191 -58 195
rect -54 193 -48 195
rect -44 193 -40 197
rect -36 193 -32 197
rect -28 193 -24 197
rect -20 193 -15 197
rect -11 193 -7 197
rect -3 193 1 197
rect 5 193 23 197
rect 27 193 31 197
rect 35 193 47 197
rect 51 193 55 197
rect 59 193 63 197
rect 67 193 71 197
rect 75 193 79 197
rect 83 195 224 197
rect 83 193 87 195
rect -54 191 87 193
rect 91 191 101 195
rect 105 191 111 195
rect 115 191 125 195
rect 129 191 135 195
rect 139 191 149 195
rect 153 191 159 195
rect 163 191 173 195
rect 177 191 184 195
rect 188 191 198 195
rect 202 193 224 195
rect 228 193 232 197
rect 236 193 240 197
rect 244 193 260 197
rect 264 193 268 197
rect 272 193 276 197
rect 280 193 284 197
rect 288 193 292 197
rect 296 195 415 197
rect 296 193 300 195
rect 202 191 300 193
rect 304 191 314 195
rect 318 191 324 195
rect 328 191 338 195
rect 342 191 348 195
rect 352 191 362 195
rect 366 191 372 195
rect 376 191 386 195
rect 390 191 397 195
rect 401 191 411 195
rect -72 190 83 191
rect 87 190 296 191
rect 300 190 415 191
rect -72 186 -68 190
rect -48 186 -44 190
rect -32 186 -28 190
rect -15 186 -11 190
rect 1 186 5 190
rect 23 186 27 190
rect 47 186 51 190
rect 63 186 67 190
rect 71 186 75 190
rect 87 186 91 190
rect 111 186 115 190
rect 135 186 139 190
rect 159 186 163 190
rect 184 186 188 190
rect 224 186 228 190
rect 240 186 244 190
rect 260 186 264 190
rect 276 186 280 190
rect 284 186 288 190
rect 300 186 304 190
rect 324 186 328 190
rect 348 186 352 190
rect 372 186 376 190
rect 397 186 401 190
rect -64 174 -54 178
rect -64 152 -60 174
rect -64 148 -47 152
rect -64 118 -60 148
rect -40 118 -36 178
rect -24 172 -20 178
rect -24 118 -20 167
rect -7 145 -3 178
rect 31 154 35 178
rect 31 149 36 154
rect -7 141 1 145
rect -7 122 -3 141
rect 12 130 17 133
rect -7 118 3 122
rect 31 118 35 149
rect 55 137 59 178
rect 55 133 72 137
rect 55 122 59 133
rect 79 125 83 178
rect 95 174 105 178
rect 119 174 129 178
rect 143 174 153 178
rect 167 174 177 178
rect 192 174 202 178
rect 95 154 99 174
rect 95 150 103 154
rect 55 118 65 122
rect 79 121 88 125
rect 79 118 83 121
rect 95 118 99 150
rect 119 145 123 174
rect 119 141 136 145
rect 119 118 123 141
rect 143 131 147 174
rect 167 170 171 174
rect 167 166 185 170
rect 143 127 160 131
rect 143 118 147 127
rect 167 118 171 166
rect 192 118 196 174
rect 232 143 236 178
rect 232 139 240 143
rect 232 122 236 139
rect 268 137 272 178
rect 268 133 285 137
rect 268 122 272 133
rect 292 125 296 178
rect 308 174 318 178
rect 332 174 342 178
rect 356 174 366 178
rect 380 174 390 178
rect 405 174 415 178
rect 308 153 312 174
rect 308 149 316 153
rect 232 118 242 122
rect 268 118 278 122
rect 292 121 301 125
rect 292 118 296 121
rect 308 118 312 149
rect 332 125 336 174
rect 356 131 360 174
rect 380 170 384 174
rect 380 166 398 170
rect 356 127 373 131
rect 332 121 349 125
rect 332 118 336 121
rect 356 118 360 127
rect 380 118 384 166
rect 405 143 409 174
rect 405 139 419 143
rect 405 118 409 139
rect -72 110 -68 114
rect -56 110 -52 114
rect -48 110 -44 114
rect -32 110 -28 114
rect -15 110 -11 114
rect 23 110 27 114
rect 47 110 51 114
rect 71 110 75 114
rect 87 110 91 114
rect 103 110 107 114
rect 111 110 115 114
rect 127 110 131 114
rect 135 110 139 114
rect 151 110 155 114
rect 159 110 163 114
rect 175 110 179 114
rect 184 110 188 114
rect 200 110 204 114
rect 224 110 228 114
rect 260 110 264 114
rect 284 110 288 114
rect 300 110 304 114
rect 316 110 320 114
rect 324 110 328 114
rect 340 110 344 114
rect 348 110 352 114
rect 364 110 368 114
rect 372 110 376 114
rect 388 110 392 114
rect 397 110 401 114
rect 413 110 417 114
rect -72 109 417 110
rect -68 105 -64 109
rect -60 105 -56 109
rect -52 107 87 109
rect -52 105 -48 107
rect -72 103 -48 105
rect -44 103 -40 107
rect -36 103 -32 107
rect -28 103 -24 107
rect -20 103 -15 107
rect -11 103 -4 107
rect 0 103 23 107
rect 27 103 31 107
rect 35 103 47 107
rect 51 103 58 107
rect 62 103 71 107
rect 75 103 79 107
rect 83 105 87 107
rect 91 105 95 109
rect 99 105 103 109
rect 107 105 111 109
rect 115 105 119 109
rect 123 105 127 109
rect 131 105 135 109
rect 139 105 143 109
rect 147 105 151 109
rect 155 105 159 109
rect 163 105 167 109
rect 171 105 175 109
rect 179 105 184 109
rect 188 105 192 109
rect 196 105 200 109
rect 204 107 300 109
rect 204 105 224 107
rect 83 103 224 105
rect 228 103 235 107
rect 239 103 260 107
rect 264 103 271 107
rect 275 103 284 107
rect 288 103 292 107
rect 296 105 300 107
rect 304 105 308 109
rect 312 105 316 109
rect 320 105 324 109
rect 328 105 332 109
rect 336 105 340 109
rect 344 105 348 109
rect 352 105 356 109
rect 360 105 364 109
rect 368 105 372 109
rect 376 105 380 109
rect 384 105 388 109
rect 392 105 397 109
rect 401 105 405 109
rect 409 105 413 109
rect 296 103 417 105
rect -72 102 417 103
<< m2contact >>
rect -24 167 -19 172
rect -36 159 -31 164
rect 36 149 41 154
rect 1 141 6 146
rect 12 125 17 130
rect 103 149 108 154
rect 240 139 245 144
rect 316 149 321 154
<< pm12contact >>
rect -15 167 -10 172
rect 0 125 5 130
rect 23 125 28 130
rect 47 125 52 130
rect 62 125 67 130
rect 102 166 107 171
rect 111 123 116 128
rect 126 132 131 137
rect 150 141 155 146
rect 174 149 179 154
rect 224 167 229 172
rect 199 158 204 163
rect 239 149 244 154
rect 260 149 265 154
rect 275 125 280 130
rect 315 166 320 171
rect 324 125 329 130
rect 339 128 344 133
rect 363 139 368 144
rect 387 149 392 154
rect 412 158 417 163
<< metal2 >>
rect -19 167 -15 171
rect -10 167 102 171
rect 107 167 224 171
rect 229 167 315 171
rect -31 158 199 162
rect 204 158 412 162
rect 34 149 36 154
rect 41 149 44 154
rect 49 149 51 154
rect 108 150 174 154
rect 244 149 249 154
rect 256 149 260 154
rect 321 150 387 154
rect 6 141 150 145
rect 245 140 363 144
rect 131 132 133 137
rect 138 132 139 137
rect 5 125 12 129
rect 17 125 23 129
rect 28 125 47 129
rect 67 125 111 129
rect 116 124 275 128
rect 280 125 324 129
rect 344 128 347 133
<< m3contact >>
rect 44 149 49 154
rect 249 149 256 154
rect 133 132 138 137
rect 347 128 352 136
<< metal3 >>
rect 49 149 249 154
rect 138 136 352 137
rect 138 132 347 136
<< labels >>
rlabel polycontact -71 167 -67 171 1 S2
rlabel polycontact -57 167 -53 171 1 RST
rlabel polycontact -31 168 -27 172 1 S1
rlabel metal1 -51 190 -51 198 1 VDD
rlabel metal1 -51 102 -51 110 1 GND
rlabel pm12contact 62 125 67 130 1 S0
rlabel pm12contact 126 132 131 137 1 REQ
rlabel metal1 415 139 419 143 7 N0
rlabel metal1 192 141 196 145 1 N1
rlabel metal1 12 130 17 133 1 T
<< end >>
