magic
tech scmos
timestamp 1732211089
<< nwell >>
rect -10 69 199 97
<< ntransistor >>
rect 2 11 4 15
rect 8 11 10 15
rect 26 11 28 15
rect 42 11 44 15
rect 50 11 52 15
rect 66 11 68 15
rect 74 11 76 15
rect 90 11 92 15
rect 96 11 98 15
rect 114 11 116 15
rect 130 11 132 15
rect 138 11 140 15
rect 154 11 156 15
rect 162 11 164 15
rect 180 11 182 15
rect 186 11 188 15
<< ptransistor >>
rect 2 75 4 83
rect 10 75 12 83
rect 26 75 28 83
rect 44 75 46 83
rect 50 75 52 83
rect 68 75 70 83
rect 74 75 76 83
rect 90 75 92 83
rect 98 75 100 83
rect 114 75 116 83
rect 132 75 134 83
rect 138 75 140 83
rect 156 75 158 83
rect 162 75 164 83
rect 178 75 180 83
rect 186 75 188 83
<< ndiffusion >>
rect 1 11 2 15
rect 4 11 8 15
rect 10 11 11 15
rect 25 11 26 15
rect 28 11 29 15
rect 41 11 42 15
rect 44 11 45 15
rect 49 11 50 15
rect 52 11 53 15
rect 65 11 66 15
rect 68 11 69 15
rect 73 11 74 15
rect 76 11 77 15
rect 89 11 90 15
rect 92 11 96 15
rect 98 11 99 15
rect 113 11 114 15
rect 116 11 117 15
rect 129 11 130 15
rect 132 11 133 15
rect 137 11 138 15
rect 140 11 141 15
rect 153 11 154 15
rect 156 11 157 15
rect 161 11 162 15
rect 164 11 165 15
rect 179 11 180 15
rect 182 11 186 15
rect 188 11 189 15
<< pdiffusion >>
rect 1 75 2 83
rect 4 75 5 83
rect 9 75 10 83
rect 12 75 13 83
rect 25 75 26 83
rect 28 75 29 83
rect 43 75 44 83
rect 46 75 50 83
rect 52 75 53 83
rect 67 75 68 83
rect 70 75 74 83
rect 76 75 77 83
rect 89 75 90 83
rect 92 75 93 83
rect 97 75 98 83
rect 100 75 101 83
rect 113 75 114 83
rect 116 75 117 83
rect 131 75 132 83
rect 134 75 138 83
rect 140 75 141 83
rect 155 75 156 83
rect 158 75 162 83
rect 164 75 165 83
rect 177 75 178 83
rect 180 75 181 83
rect 185 75 186 83
rect 188 75 189 83
<< ndcontact >>
rect -3 11 1 15
rect 11 11 15 15
rect 21 11 25 15
rect 29 11 33 15
rect 37 11 41 15
rect 45 11 49 15
rect 53 11 57 15
rect 61 11 65 15
rect 69 11 73 15
rect 77 11 81 15
rect 85 11 89 15
rect 99 11 103 15
rect 109 11 113 15
rect 117 11 121 15
rect 125 11 129 15
rect 133 11 137 15
rect 141 11 145 15
rect 149 11 153 15
rect 157 11 161 15
rect 165 11 169 15
rect 175 11 179 15
rect 189 11 193 15
<< pdcontact >>
rect -3 75 1 83
rect 5 75 9 83
rect 13 75 17 83
rect 21 75 25 83
rect 29 75 33 83
rect 39 75 43 83
rect 53 75 57 83
rect 63 75 67 83
rect 77 75 81 83
rect 85 75 89 83
rect 93 75 97 83
rect 101 75 105 83
rect 109 75 113 83
rect 117 75 121 83
rect 127 75 131 83
rect 141 75 145 83
rect 151 75 155 83
rect 165 75 169 83
rect 173 75 177 83
rect 181 75 185 83
rect 189 75 193 83
<< psubstratepcontact >>
rect -3 0 1 4
rect 8 0 12 4
rect 21 0 25 4
rect 29 0 33 4
rect 37 0 41 4
rect 45 0 49 4
rect 53 0 57 4
rect 61 0 65 4
rect 69 0 73 4
rect 77 0 81 4
rect 85 0 89 4
rect 96 0 100 4
rect 109 0 113 4
rect 117 0 121 4
rect 125 0 129 4
rect 133 0 137 4
rect 141 0 145 4
rect 149 0 153 4
rect 157 0 161 4
rect 165 0 169 4
rect 178 0 182 4
rect 189 0 193 4
<< nsubstratencontact >>
rect -3 90 1 94
rect 5 90 9 94
rect 13 90 17 94
rect 21 90 25 94
rect 29 90 33 94
rect 39 90 43 94
rect 53 90 57 94
rect 63 90 67 94
rect 77 90 81 94
rect 85 90 89 94
rect 93 90 97 94
rect 101 90 105 94
rect 109 90 113 94
rect 117 90 121 94
rect 127 90 131 94
rect 141 90 145 94
rect 151 90 155 94
rect 165 90 169 94
rect 173 90 177 94
rect 181 90 185 94
rect 189 90 193 94
<< polysilicon >>
rect 2 83 4 86
rect 10 83 12 86
rect 26 83 28 86
rect 44 83 46 86
rect 50 83 52 86
rect 68 83 70 86
rect 74 83 76 86
rect 90 83 92 86
rect 98 83 100 86
rect 114 83 116 86
rect 132 83 134 86
rect 138 83 140 86
rect 156 83 158 86
rect 162 83 164 86
rect 178 83 180 86
rect 186 83 188 86
rect 2 15 4 75
rect 10 23 12 75
rect 26 49 28 75
rect 44 50 46 75
rect 25 45 28 49
rect 8 21 12 23
rect 8 15 10 21
rect 26 15 28 45
rect 42 48 46 50
rect 42 15 44 48
rect 50 15 52 75
rect 68 44 70 75
rect 66 42 70 44
rect 66 15 68 42
rect 74 15 76 75
rect 90 15 92 75
rect 98 23 100 75
rect 114 42 116 75
rect 132 50 134 75
rect 113 38 116 42
rect 96 21 100 23
rect 96 15 98 21
rect 114 15 116 38
rect 130 48 134 50
rect 130 15 132 48
rect 138 15 140 75
rect 156 44 158 75
rect 154 42 158 44
rect 154 15 156 42
rect 162 15 164 75
rect 178 27 180 75
rect 178 25 182 27
rect 180 15 182 25
rect 186 15 188 75
rect 2 8 4 11
rect 8 8 10 11
rect 26 8 28 11
rect 42 8 44 11
rect 50 8 52 11
rect 66 8 68 11
rect 74 8 76 11
rect 90 8 92 11
rect 96 8 98 11
rect 114 8 116 11
rect 130 8 132 11
rect 138 8 140 11
rect 154 8 156 11
rect 162 8 164 11
rect 180 8 182 11
rect 186 8 188 11
<< polycontact >>
rect 21 45 25 49
rect 38 26 42 30
rect 52 26 56 30
rect 109 38 113 42
rect 126 26 130 30
rect 140 26 144 30
<< metal1 >>
rect -3 94 193 95
rect 1 90 5 94
rect 9 90 13 94
rect 17 90 21 94
rect 25 90 29 94
rect 33 90 39 94
rect 43 90 53 94
rect 57 90 63 94
rect 67 90 77 94
rect 81 90 85 94
rect 89 90 93 94
rect 97 90 101 94
rect 105 90 109 94
rect 113 90 117 94
rect 121 90 127 94
rect 131 90 141 94
rect 145 90 151 94
rect 155 90 165 94
rect 169 90 173 94
rect 177 90 181 94
rect 185 90 189 94
rect -3 87 193 90
rect -3 83 1 87
rect 13 83 17 87
rect 21 83 25 87
rect 53 83 57 87
rect 77 83 81 87
rect 5 32 9 75
rect 21 32 25 45
rect 5 27 13 32
rect 18 27 25 32
rect 29 30 33 75
rect 85 83 89 87
rect 101 83 105 87
rect 109 83 113 87
rect 141 83 145 87
rect 165 83 169 87
rect 39 55 43 75
rect 37 51 43 55
rect 63 53 67 75
rect 37 44 41 51
rect 61 49 67 53
rect 41 40 49 44
rect 13 20 17 27
rect 11 17 17 20
rect 29 26 38 30
rect 11 15 15 17
rect 29 15 33 26
rect 45 15 49 40
rect 61 30 65 49
rect 93 33 97 75
rect 109 33 113 38
rect 56 26 73 30
rect 93 28 101 33
rect 106 29 113 33
rect 117 30 121 75
rect 173 83 177 87
rect 189 83 193 87
rect 127 55 131 75
rect 125 51 131 55
rect 151 53 155 75
rect 125 44 129 51
rect 149 49 155 53
rect 124 40 137 44
rect 124 39 129 40
rect 69 15 73 26
rect 101 20 105 28
rect 99 17 105 20
rect 117 26 126 30
rect 99 15 103 17
rect 117 15 121 26
rect 133 15 137 40
rect 149 30 153 49
rect 181 41 185 75
rect 173 36 185 41
rect 173 33 177 36
rect 144 26 161 30
rect 168 28 177 33
rect 157 15 161 26
rect 173 22 177 28
rect 173 18 179 22
rect 175 15 179 18
rect -3 7 1 11
rect 21 7 25 11
rect 37 7 41 11
rect 53 7 57 11
rect 61 7 65 11
rect 77 7 81 11
rect 85 7 89 11
rect 109 7 113 11
rect 125 7 129 11
rect 141 7 145 11
rect 149 7 153 11
rect 165 7 169 11
rect 189 7 193 11
rect -3 4 193 7
rect 1 0 8 4
rect 12 0 21 4
rect 25 0 29 4
rect 33 0 37 4
rect 41 0 45 4
rect 49 0 53 4
rect 57 0 61 4
rect 65 0 69 4
rect 73 0 77 4
rect 81 0 85 4
rect 89 0 96 4
rect 100 0 109 4
rect 113 0 117 4
rect 121 0 125 4
rect 129 0 133 4
rect 137 0 141 4
rect 145 0 149 4
rect 153 0 157 4
rect 161 0 165 4
rect 169 0 178 4
rect 182 0 189 4
rect -3 -1 193 0
<< m2contact >>
rect 13 27 18 32
rect 101 28 106 33
<< pm12contact >>
rect 12 62 17 67
rect 76 62 81 67
rect -3 18 2 23
rect 100 62 105 67
rect 164 62 169 67
rect 173 54 178 59
rect 61 18 66 23
rect 85 18 90 23
rect 188 45 193 50
rect 149 18 154 23
<< ndm12contact >>
rect 36 39 41 44
<< metal2 >>
rect 17 62 76 67
rect 105 62 164 67
rect 13 54 173 58
rect 13 32 17 54
rect 101 45 188 49
rect 41 39 83 44
rect 79 23 83 39
rect 101 33 105 45
rect 2 18 61 23
rect 79 18 85 23
rect 90 18 149 23
<< labels >>
rlabel nwell -3 87 17 95 1 VDD
rlabel metal2 17 65 17 67 1 B
rlabel metal2 -3 21 -3 23 1 A
rlabel metal1 4 2 4 2 1 GND
rlabel metal2 105 65 105 67 1 C
rlabel metal1 127 42 127 42 1 Sum
rlabel metal1 171 30 171 30 1 Cout
<< end >>
