module not_gate_32 (
  output[31:0] result,
  input [31:0] a
);

  not not_0(result[0], a[0]);
  not not_1(result[1], a[1]);
  not not_2(result[2], a[2]);
  not not_3(result[3], a[3]);
  not not_4(result[4], a[4]);
  not not_5(result[5], a[5]);
  not not_6(result[6], a[6]);
  not not_7(result[7], a[7]);
  not not_8(result[8], a[8]);
  not not_9(result[9], a[9]);
  not not_10(result[10], a[10]);
  not not_11(result[11], a[11]);
  not not_12(result[12], a[12]);
  not not_13(result[13], a[13]);
  not not_14(result[14], a[14]);
  not not_15(result[15], a[15]);
  not not_16(result[16], a[16]);
  not not_17(result[17], a[17]);
  not not_18(result[18], a[18]);
  not not_19(result[19], a[19]);
  not not_20(result[20], a[20]);
  not not_21(result[21], a[21]);
  not not_22(result[22], a[22]);
  not not_23(result[23], a[23]);
  not not_24(result[24], a[24]);
  not not_25(result[25], a[25]);
  not not_26(result[26], a[26]);
  not not_27(result[27], a[27]);
  not not_28(result[28], a[28]);
  not not_29(result[29], a[29]);
  not not_30(result[30], a[30]);
  not not_31(result[31], a[31]);

endmodule
