module CLA_32bit_2level();









endmodule 