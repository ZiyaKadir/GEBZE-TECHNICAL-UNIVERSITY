magic
tech scmos
timestamp 1734635707
<< nwell >>
rect -70 29 218 61
<< ntransistor >>
rect -59 -38 -57 -34
rect -37 -36 -35 -32
rect -5 -38 -3 -34
rect 1 -38 3 -34
rect 9 -38 11 -34
rect 45 -38 47 -34
rect 53 -38 55 -34
rect 59 -38 61 -34
rect 82 -38 84 -34
rect 107 -36 109 -32
rect 140 -38 142 -34
rect 146 -38 148 -34
rect 154 -38 156 -34
rect 189 -38 191 -34
rect 197 -38 199 -34
rect 203 -38 205 -34
<< ptransistor >>
rect -59 35 -57 43
rect -37 35 -35 43
rect -5 35 -3 43
rect 3 35 5 43
rect 11 35 13 43
rect 43 35 45 43
rect 51 35 53 43
rect 59 35 61 43
rect 82 35 84 43
rect 107 35 109 43
rect 140 35 142 43
rect 148 35 150 43
rect 156 35 158 43
rect 187 35 189 43
rect 195 35 197 43
rect 203 35 205 43
<< ndiffusion >>
rect -60 -38 -59 -34
rect -57 -38 -56 -34
rect -38 -36 -37 -32
rect -35 -36 -34 -32
rect -6 -38 -5 -34
rect -3 -38 1 -34
rect 3 -38 4 -34
rect 8 -38 9 -34
rect 11 -38 12 -34
rect 44 -38 45 -34
rect 47 -38 48 -34
rect 52 -38 53 -34
rect 55 -38 59 -34
rect 61 -38 62 -34
rect 81 -38 82 -34
rect 84 -38 85 -34
rect 106 -36 107 -32
rect 109 -36 110 -32
rect 139 -38 140 -34
rect 142 -38 146 -34
rect 148 -38 149 -34
rect 153 -38 154 -34
rect 156 -38 157 -34
rect 188 -38 189 -34
rect 191 -38 192 -34
rect 196 -38 197 -34
rect 199 -38 203 -34
rect 205 -38 206 -34
<< pdiffusion >>
rect -60 35 -59 43
rect -57 35 -56 43
rect -38 35 -37 43
rect -35 35 -34 43
rect -6 35 -5 43
rect -3 35 -2 43
rect 2 35 3 43
rect 5 35 6 43
rect 10 35 11 43
rect 13 35 14 43
rect 42 35 43 43
rect 45 35 46 43
rect 50 35 51 43
rect 53 35 54 43
rect 58 35 59 43
rect 61 35 62 43
rect 81 35 82 43
rect 84 35 85 43
rect 106 35 107 43
rect 109 35 110 43
rect 139 35 140 43
rect 142 35 143 43
rect 147 35 148 43
rect 150 35 151 43
rect 155 35 156 43
rect 158 35 159 43
rect 186 35 187 43
rect 189 35 190 43
rect 194 35 195 43
rect 197 35 198 43
rect 202 35 203 43
rect 205 35 206 43
<< ndcontact >>
rect -64 -38 -60 -34
rect -56 -38 -52 -34
rect -42 -36 -38 -32
rect -34 -36 -30 -32
rect -10 -38 -6 -34
rect 4 -38 8 -34
rect 12 -38 16 -34
rect 40 -38 44 -34
rect 48 -38 52 -34
rect 62 -38 66 -34
rect 77 -38 81 -34
rect 85 -38 89 -34
rect 102 -36 106 -32
rect 110 -36 114 -32
rect 135 -38 139 -34
rect 149 -38 153 -34
rect 157 -38 161 -34
rect 184 -38 188 -34
rect 192 -38 196 -34
rect 206 -38 210 -34
<< pdcontact >>
rect -64 35 -60 43
rect -56 35 -52 43
rect -42 35 -38 43
rect -34 35 -30 43
rect -10 35 -6 43
rect -2 35 2 43
rect 6 35 10 43
rect 14 35 18 43
rect 38 35 42 43
rect 46 35 50 43
rect 54 35 58 43
rect 62 35 66 43
rect 77 35 81 43
rect 85 35 89 43
rect 102 35 106 43
rect 110 35 114 43
rect 135 35 139 43
rect 143 35 147 43
rect 151 35 155 43
rect 159 35 163 43
rect 182 35 186 43
rect 190 35 194 43
rect 198 35 202 43
rect 206 35 210 43
<< psubstratepcontact >>
rect -64 -48 -60 -44
rect -56 -48 -52 -44
rect -42 -48 -38 -44
rect -34 -48 -30 -44
rect -10 -48 -6 -44
rect 4 -48 8 -44
rect 12 -48 16 -44
rect 40 -48 44 -44
rect 48 -48 52 -44
rect 62 -48 66 -44
rect 77 -48 81 -44
rect 85 -48 89 -44
rect 102 -48 106 -44
rect 110 -48 114 -44
rect 135 -48 139 -44
rect 149 -48 153 -44
rect 157 -48 161 -44
rect 184 -48 188 -44
rect 192 -48 196 -44
rect 206 -48 210 -44
<< nsubstratencontact >>
rect -64 49 -60 53
rect -56 49 -52 53
rect -42 49 -38 53
rect -34 49 -30 53
rect -10 49 -6 53
rect -2 49 2 53
rect 6 49 10 53
rect 14 49 18 53
rect 38 49 42 53
rect 46 49 50 53
rect 54 49 58 53
rect 62 49 66 53
rect 102 49 106 53
rect 110 49 114 53
rect 135 49 139 53
rect 143 49 147 53
rect 151 49 155 53
rect 159 49 163 53
rect 182 49 186 53
rect 190 49 194 53
rect 198 49 202 53
rect 206 49 210 53
<< polysilicon >>
rect -59 43 -57 46
rect -37 43 -35 46
rect -5 43 -3 46
rect 3 43 5 46
rect 11 43 13 46
rect 43 43 45 46
rect 51 43 53 46
rect 59 43 61 46
rect 82 43 84 46
rect 107 43 109 46
rect 140 43 142 46
rect 148 43 150 46
rect 156 43 158 46
rect 187 43 189 46
rect 195 43 197 46
rect 203 43 205 46
rect -59 -34 -57 35
rect -37 17 -35 35
rect -5 17 -3 35
rect 3 24 5 35
rect -37 13 -34 17
rect -37 -32 -35 13
rect -5 -34 -3 13
rect 3 9 5 19
rect 0 7 5 9
rect 0 -31 2 7
rect 11 -13 13 35
rect 43 1 45 35
rect 51 11 53 35
rect 59 24 61 35
rect 43 -1 47 1
rect 9 -15 13 -13
rect 0 -33 3 -31
rect 1 -34 3 -33
rect 9 -34 11 -15
rect 45 -34 47 -1
rect 51 0 53 6
rect 51 -2 55 0
rect 53 -34 55 -2
rect 59 -34 61 19
rect 82 -34 84 35
rect 107 -32 109 35
rect 140 -6 142 35
rect 148 24 150 35
rect 148 9 150 19
rect 141 -10 142 -6
rect -59 -41 -57 -38
rect -37 -39 -35 -36
rect 140 -34 142 -10
rect 145 7 150 9
rect 145 -31 147 7
rect 156 -13 158 35
rect 187 1 189 35
rect 195 11 197 35
rect 203 24 205 35
rect 187 -1 191 1
rect 154 -15 158 -13
rect 145 -33 148 -31
rect 146 -34 148 -33
rect 154 -34 156 -15
rect 189 -34 191 -1
rect 195 0 197 6
rect 195 -2 199 0
rect 197 -34 199 -2
rect 203 -34 205 19
rect -5 -41 -3 -38
rect 1 -41 3 -38
rect 9 -41 11 -38
rect 45 -41 47 -38
rect 53 -41 55 -38
rect 59 -41 61 -38
rect 82 -41 84 -38
rect 107 -39 109 -36
rect 140 -41 142 -38
rect 146 -41 148 -38
rect 154 -41 156 -38
rect 189 -41 191 -38
rect 197 -41 199 -38
rect 203 -41 205 -38
<< polycontact >>
rect -63 -6 -59 -2
rect -34 13 -30 17
rect -7 13 -3 17
rect 78 20 82 24
rect 41 -21 45 -17
rect 137 -10 141 -6
rect 185 -21 189 -17
<< metal1 >>
rect -66 53 212 55
rect -66 49 -64 53
rect -60 49 -56 53
rect -52 49 -42 53
rect -38 49 -34 53
rect -30 49 -10 53
rect -6 49 -2 53
rect 2 49 6 53
rect 10 49 14 53
rect 18 49 38 53
rect 42 49 46 53
rect 50 49 54 53
rect 58 49 62 53
rect 66 49 102 53
rect 106 49 110 53
rect 114 49 135 53
rect 139 49 143 53
rect 147 49 151 53
rect 155 49 159 53
rect 163 49 182 53
rect 186 49 190 53
rect 194 49 198 53
rect 202 49 206 53
rect 210 49 212 53
rect -66 47 212 49
rect -64 43 -60 47
rect -34 43 -30 47
rect -2 43 2 47
rect 54 43 58 47
rect 77 43 81 47
rect 110 43 114 47
rect 143 43 147 47
rect 198 43 202 47
rect -56 25 -52 35
rect -56 -34 -52 20
rect -42 11 -38 35
rect -10 31 -6 35
rect 6 31 10 35
rect -10 27 10 31
rect -30 13 -7 17
rect -41 6 -38 11
rect -42 -32 -38 6
rect 14 -17 18 35
rect 38 -4 42 35
rect 46 31 50 35
rect 62 31 66 35
rect 46 27 66 31
rect 62 20 78 24
rect 43 -9 52 -5
rect 4 -21 41 -17
rect 4 -34 8 -21
rect 48 -34 52 -9
rect 85 -34 89 35
rect 102 11 106 35
rect 135 31 139 35
rect 151 31 155 35
rect 135 27 155 31
rect 103 6 106 11
rect -64 -42 -60 -38
rect -34 -42 -30 -36
rect -10 -42 -6 -38
rect 12 -42 16 -38
rect 40 -42 44 -38
rect 62 -42 66 -38
rect 102 -32 106 6
rect 114 -10 137 -6
rect 159 -17 163 35
rect 182 -4 186 35
rect 190 31 194 35
rect 206 31 210 35
rect 190 27 210 31
rect 187 -9 196 -5
rect 149 -21 185 -17
rect 149 -34 153 -21
rect 192 -34 196 -9
rect 77 -42 81 -38
rect 110 -42 114 -36
rect 135 -42 139 -38
rect 157 -42 161 -38
rect 184 -42 188 -38
rect 206 -42 210 -38
rect -66 -44 212 -42
rect -66 -48 -64 -44
rect -60 -48 -56 -44
rect -52 -48 -42 -44
rect -38 -48 -34 -44
rect -30 -48 -10 -44
rect -6 -48 4 -44
rect 8 -48 12 -44
rect 16 -48 40 -44
rect 44 -48 48 -44
rect 52 -48 62 -44
rect 66 -48 77 -44
rect 81 -48 85 -44
rect 89 -48 102 -44
rect 106 -48 110 -44
rect 114 -48 135 -44
rect 139 -48 149 -44
rect 153 -48 157 -44
rect 161 -48 184 -44
rect 188 -48 192 -44
rect 196 -48 206 -44
rect 210 -48 212 -44
rect -66 -50 212 -48
<< m2contact >>
rect -56 20 -51 25
rect -46 6 -41 11
rect 38 -9 43 -4
rect 89 20 94 25
rect 98 6 103 11
rect 182 -9 187 -4
<< pm12contact >>
rect 1 19 6 24
rect 6 -9 11 -4
rect 57 19 62 24
rect 49 6 54 11
rect 146 19 151 24
rect 109 -10 114 -5
rect 151 -9 156 -4
rect 201 19 206 24
rect 193 6 198 11
<< metal2 >>
rect -51 20 1 24
rect 6 20 57 24
rect 94 20 146 24
rect 151 20 201 24
rect -41 6 49 10
rect 103 6 193 10
rect 11 -9 38 -5
rect 43 -9 109 -5
rect 156 -9 182 -5
<< labels >>
rlabel pm12contact 154 -7 154 -7 1 Q
rlabel polycontact 187 -19 187 -19 1 notQ
rlabel polycontact -5 15 -5 15 1 D
rlabel polycontact -61 -4 -61 -4 1 CLK
rlabel metal1 28 51 28 51 1 VDD
rlabel metal1 26 -46 26 -46 1 GND
<< end >>
