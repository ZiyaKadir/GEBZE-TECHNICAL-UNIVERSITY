module nor_gate_32 (
output [31:0]result, 
input [31:0]a,
input [31:0]b
);
	
	
	nor nor_0(result[0],a[0],b[0]);
	nor nor_1(result[1],a[1],b[1]);
	nor nor_2(result[2],a[2],b[2]);
	nor nor_3(result[3],a[3],b[3]);
	nor nor_4(result[4],a[4],b[4]);
	nor nor_5(result[5],a[5],b[5]);
	nor nor_6(result[6],a[6],b[6]);
	nor nor_7(result[7],a[7],b[7]);
	nor nor_8(result[8],a[8],b[8]);
	nor nor_9(result[9],a[9],b[9]);
	nor nor_10(result[10],a[10],b[10]);
	nor nor_11(result[11],a[11],b[11]);
	nor nor_12(result[12],a[12],b[12]);
	nor nor_13(result[13],a[13],b[13]);
	nor nor_14(result[14],a[14],b[14]);
	nor nor_15(result[15],a[15],b[15]);
	nor nor_16(result[16],a[16],b[16]);
	nor nor_17(result[17],a[17],b[17]);
	nor nor_18(result[18],a[18],b[18]);
	nor nor_19(result[19],a[19],b[19]);
	nor nor_20(result[20],a[20],b[20]);
	nor nor_21(result[21],a[21],b[21]);
	nor nor_22(result[22],a[22],b[22]);
	nor nor_23(result[23],a[23],b[23]);
	nor nor_24(result[24],a[24],b[24]);
	nor nor_25(result[25],a[25],b[25]);
	nor nor_26(result[26],a[26],b[26]);
	nor nor_27(result[27],a[27],b[27]);
	nor nor_28(result[28],a[28],b[28]);
	nor nor_29(result[29],a[29],b[29]);
	nor nor_30(result[30],a[30],b[30]);
	nor nor_31(result[31],a[31],b[31]);

	
endmodule 