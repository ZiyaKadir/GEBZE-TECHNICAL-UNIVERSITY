module _4or(

	input a,
	input b,
	input c,
	input d,
	
	output out
);

	or res_or(out,a,b,c,d);

endmodule 