magic
tech scmos
timestamp 1730394342
<< nwell >>
rect -16 20 14 48
<< ntransistor >>
rect -5 -39 -3 -35
rect 3 -39 5 -35
<< ptransistor >>
rect -5 26 -3 34
rect 1 26 3 34
<< ndiffusion >>
rect -6 -39 -5 -35
rect -3 -39 -2 -35
rect 2 -39 3 -35
rect 5 -39 6 -35
<< pdiffusion >>
rect -6 26 -5 34
rect -3 26 1 34
rect 3 26 4 34
<< ndcontact >>
rect -10 -39 -6 -35
rect -2 -39 2 -35
rect 6 -39 10 -35
<< pdcontact >>
rect -10 26 -6 34
rect 4 26 8 34
<< psubstratepcontact >>
rect -10 -48 -6 -44
rect -2 -48 2 -44
rect 6 -48 10 -44
<< nsubstratencontact >>
rect -10 39 -6 43
rect 4 39 8 43
<< polysilicon >>
rect -5 34 -3 37
rect 1 34 3 37
rect -5 -35 -3 26
rect 1 -6 3 26
rect 1 -8 5 -6
rect 3 -35 5 -8
rect -5 -42 -3 -39
rect 3 -42 5 -39
<< polycontact >>
rect -9 -3 -5 1
rect 5 -27 9 -23
<< metal1 >>
rect -10 43 8 46
rect -6 39 4 43
rect -10 38 8 39
rect -10 34 -6 38
rect 4 3 8 26
rect 4 -1 10 3
rect 6 -4 10 -1
rect 6 -8 14 -4
rect 6 -12 10 -8
rect -2 -16 10 -12
rect -2 -35 2 -16
rect -10 -43 -6 -39
rect 6 -43 10 -39
rect -10 -44 10 -43
rect -6 -48 -2 -44
rect 2 -48 6 -44
rect -10 -51 10 -48
<< labels >>
rlabel polycontact -9 -3 -5 1 1 A
rlabel polycontact 5 -27 9 -23 1 B
rlabel metal1 10 -8 14 -4 7 Y
rlabel metal1 -10 -51 10 -43 1 GND
rlabel nwell -10 38 8 46 1 VDD
<< end >>
