* SPICE3 file created from HW_1_NAND.ext - technology: scmos

.option scale=0.12u
.include tsmc_cmos025

.model nfet NMOS
.model pfet PMOS

Vdd VDD 0 2.5V
Vina A 0 PULSE(0 2.5 0ns 10ns 10ns 20ns 40ns)
Vinb B 0 PULSE(0 2.5 0ns 20ns 20ns 40ns 80ns)
CL Y 0 1fF
.TRAN 1ns 400ns

M1000 Y A VDD VDD pfet w=8 l=2
+  ad=24p pd=14u as=40p ps=26u
M1001 VDD B Y VDD pfet w=8 l=2
+  ad=40p pd=26u as=24p ps=14u
M1002 Y B a_n3_n42# Gnd nfet w=4 l=2
+  ad=20p pd=18u as=8p ps=8u
M1003 a_n3_n42# A GND Gnd nfet w=4 l=2
+  ad=8p pd=8u as=20p ps=18u
C0 A B 0.351754f
C1 B Y 0.121112f
C2 A Y 0.048377f
C3 B VDD 0.042197f
C4 A VDD 0.042197f
C5 VDD Y 0.248945f
C6 GND Y 0.011598f
C7 GND 0 0.167227f 
C8 Y 0 0.417784f 
C9 B 0 0.514983f 
C10 A 0 0.503383f 
C11 VDD 0 0.976475f 
