magic
tech scmos
timestamp 1736872262
<< nwell >>
rect -55 53 193 81
<< ntransistor >>
rect -44 -5 -42 -1
rect -36 -5 -34 -1
rect -20 -5 -18 -1
rect -4 -5 -2 -1
rect 13 -5 15 -1
rect 19 -5 21 -1
rect 37 -5 39 -1
rect 43 -5 45 -1
rect 61 -5 63 -1
rect 77 -5 79 -1
rect 85 -5 87 -1
rect 101 -5 103 -1
rect 109 -5 111 -1
rect 125 -5 127 -1
rect 133 -5 135 -1
rect 149 -5 151 -1
rect 157 -5 159 -1
rect 174 -5 176 -1
rect 182 -5 184 -1
<< ptransistor >>
rect -44 59 -42 67
rect -38 59 -36 67
rect -20 59 -18 67
rect -4 59 -2 67
rect 13 59 15 67
rect 21 59 23 67
rect 37 59 39 67
rect 45 59 47 67
rect 61 59 63 67
rect 77 59 79 67
rect 83 59 85 67
rect 101 59 103 67
rect 107 59 109 67
rect 125 59 127 67
rect 131 59 133 67
rect 149 59 151 67
rect 155 59 157 67
rect 174 59 176 67
rect 180 59 182 67
<< ndiffusion >>
rect -45 -5 -44 -1
rect -42 -5 -41 -1
rect -37 -5 -36 -1
rect -34 -5 -33 -1
rect -21 -5 -20 -1
rect -18 -5 -17 -1
rect -5 -5 -4 -1
rect -2 -5 -1 -1
rect 12 -5 13 -1
rect 15 -5 19 -1
rect 21 -5 22 -1
rect 36 -5 37 -1
rect 39 -5 43 -1
rect 45 -5 46 -1
rect 60 -5 61 -1
rect 63 -5 64 -1
rect 76 -5 77 -1
rect 79 -5 80 -1
rect 84 -5 85 -1
rect 87 -5 88 -1
rect 100 -5 101 -1
rect 103 -5 104 -1
rect 108 -5 109 -1
rect 111 -5 112 -1
rect 124 -5 125 -1
rect 127 -5 128 -1
rect 132 -5 133 -1
rect 135 -5 136 -1
rect 148 -5 149 -1
rect 151 -5 152 -1
rect 156 -5 157 -1
rect 159 -5 160 -1
rect 173 -5 174 -1
rect 176 -5 177 -1
rect 181 -5 182 -1
rect 184 -5 185 -1
<< pdiffusion >>
rect -45 59 -44 67
rect -42 59 -38 67
rect -36 59 -35 67
rect -21 59 -20 67
rect -18 59 -17 67
rect -5 59 -4 67
rect -2 59 -1 67
rect 12 59 13 67
rect 15 59 16 67
rect 20 59 21 67
rect 23 59 24 67
rect 36 59 37 67
rect 39 59 40 67
rect 44 59 45 67
rect 47 59 48 67
rect 60 59 61 67
rect 63 59 64 67
rect 76 59 77 67
rect 79 59 83 67
rect 85 59 86 67
rect 100 59 101 67
rect 103 59 107 67
rect 109 59 110 67
rect 124 59 125 67
rect 127 59 131 67
rect 133 59 134 67
rect 148 59 149 67
rect 151 59 155 67
rect 157 59 158 67
rect 173 59 174 67
rect 176 59 180 67
rect 182 59 183 67
<< ndcontact >>
rect -49 -5 -45 -1
rect -41 -5 -37 -1
rect -33 -5 -29 -1
rect -25 -5 -21 -1
rect -17 -5 -13 -1
rect -9 -5 -5 -1
rect -1 -5 3 -1
rect 8 -5 12 -1
rect 22 -5 26 -1
rect 32 -5 36 -1
rect 46 -5 50 -1
rect 56 -5 60 -1
rect 64 -5 68 -1
rect 72 -5 76 -1
rect 80 -5 84 -1
rect 88 -5 92 -1
rect 96 -5 100 -1
rect 104 -5 108 -1
rect 112 -5 116 -1
rect 120 -5 124 -1
rect 128 -5 132 -1
rect 136 -5 140 -1
rect 144 -5 148 -1
rect 152 -5 156 -1
rect 160 -5 164 -1
rect 169 -5 173 -1
rect 177 -5 181 -1
rect 185 -5 189 -1
<< pdcontact >>
rect -49 59 -45 67
rect -35 59 -31 67
rect -25 59 -21 67
rect -17 59 -13 67
rect -9 59 -5 67
rect -1 59 3 67
rect 8 59 12 67
rect 16 59 20 67
rect 24 59 28 67
rect 32 59 36 67
rect 40 59 44 67
rect 48 59 52 67
rect 56 59 60 67
rect 64 59 68 67
rect 72 59 76 67
rect 86 59 90 67
rect 96 59 100 67
rect 110 59 114 67
rect 120 59 124 67
rect 134 59 138 67
rect 144 59 148 67
rect 158 59 162 67
rect 169 59 173 67
rect 183 59 187 67
<< psubstratepcontact >>
rect -49 -14 -45 -10
rect -41 -14 -37 -10
rect -33 -14 -29 -10
rect -25 -16 -21 -12
rect -17 -16 -13 -12
rect -9 -16 -5 -12
rect -1 -16 3 -12
rect 8 -16 12 -12
rect 19 -16 23 -12
rect 32 -16 36 -12
rect 43 -16 47 -12
rect 56 -16 60 -12
rect 64 -16 68 -12
rect 72 -14 76 -10
rect 80 -14 84 -10
rect 88 -14 92 -10
rect 96 -14 100 -10
rect 104 -14 108 -10
rect 112 -14 116 -10
rect 120 -14 124 -10
rect 128 -14 132 -10
rect 136 -14 140 -10
rect 144 -14 148 -10
rect 152 -14 156 -10
rect 160 -14 164 -10
rect 169 -14 173 -10
rect 177 -14 181 -10
rect 185 -14 189 -10
<< nsubstratencontact >>
rect -49 72 -45 76
rect -35 72 -31 76
rect -25 74 -21 78
rect -17 74 -13 78
rect -9 74 -5 78
rect -1 74 3 78
rect 8 74 12 78
rect 16 74 20 78
rect 24 74 28 78
rect 32 74 36 78
rect 40 74 44 78
rect 48 74 52 78
rect 56 74 60 78
rect 64 74 68 78
rect 72 72 76 76
rect 86 72 90 76
rect 96 72 100 76
rect 110 72 114 76
rect 120 72 124 76
rect 134 72 138 76
rect 144 72 148 76
rect 158 72 162 76
rect 169 72 173 76
rect 183 72 187 76
<< polysilicon >>
rect -44 67 -42 70
rect -38 67 -36 70
rect -20 67 -18 70
rect -4 67 -2 70
rect 13 67 15 70
rect 21 67 23 70
rect 37 67 39 70
rect 45 67 47 70
rect 61 67 63 70
rect 77 67 79 70
rect 83 67 85 70
rect 101 67 103 70
rect 107 67 109 70
rect 125 67 127 70
rect 131 67 133 70
rect 149 67 151 70
rect 155 67 157 70
rect 174 67 176 70
rect 180 67 182 70
rect -44 -1 -42 59
rect -38 58 -36 59
rect -38 56 -34 58
rect -36 -1 -34 56
rect -20 -1 -18 59
rect -4 -1 -2 59
rect 13 -1 15 59
rect 21 3 23 59
rect 19 1 23 3
rect 19 -1 21 1
rect 37 -1 39 59
rect 45 3 47 59
rect 43 1 47 3
rect 43 -1 45 1
rect 61 -1 63 59
rect 77 -1 79 59
rect 83 58 85 59
rect 83 56 87 58
rect 85 -1 87 56
rect 101 -1 103 59
rect 107 58 109 59
rect 107 56 111 58
rect 109 -1 111 56
rect 125 -1 127 59
rect 131 58 133 59
rect 131 56 135 58
rect 133 -1 135 56
rect 149 -1 151 59
rect 155 58 157 59
rect 155 56 159 58
rect 157 -1 159 56
rect 174 -1 176 59
rect 180 58 182 59
rect 180 56 184 58
rect 182 -1 184 56
rect -44 -8 -42 -5
rect -36 -8 -34 -5
rect -20 -8 -18 -5
rect -4 -8 -2 -5
rect 13 -8 15 -5
rect 19 -8 21 -5
rect 37 -8 39 -5
rect 43 -8 45 -5
rect 61 -8 63 -5
rect 77 -8 79 -5
rect 85 -8 87 -5
rect 101 -8 103 -5
rect 109 -8 111 -5
rect 125 -8 127 -5
rect 133 -8 135 -5
rect 149 -8 151 -5
rect 157 -8 159 -5
rect 174 -8 176 -5
rect 182 -8 184 -5
<< polycontact >>
rect -48 48 -44 52
rect -34 48 -30 52
rect -24 29 -20 33
rect -8 49 -4 53
rect 23 6 27 10
rect 33 6 37 10
rect 57 14 61 18
rect 73 2 77 6
rect 121 12 125 16
rect 111 4 115 8
rect 145 8 149 12
rect 170 47 174 51
<< metal1 >>
rect -49 78 187 79
rect -49 76 -25 78
rect -45 72 -35 76
rect -31 74 -25 76
rect -21 74 -17 78
rect -13 74 -9 78
rect -5 74 -1 78
rect 3 74 8 78
rect 12 74 16 78
rect 20 74 24 78
rect 28 74 32 78
rect 36 74 40 78
rect 44 74 48 78
rect 52 74 56 78
rect 60 74 64 78
rect 68 76 187 78
rect 68 74 72 76
rect -31 72 72 74
rect 76 72 86 76
rect 90 72 96 76
rect 100 72 110 76
rect 114 72 120 76
rect 124 72 134 76
rect 138 72 144 76
rect 148 72 158 76
rect 162 72 169 76
rect 173 72 183 76
rect -49 71 68 72
rect 72 71 187 72
rect -49 67 -45 71
rect -25 67 -21 71
rect -9 67 -5 71
rect 8 67 12 71
rect 24 67 28 71
rect 32 67 36 71
rect 48 67 52 71
rect 56 67 60 71
rect 72 67 76 71
rect 96 67 100 71
rect 120 67 124 71
rect 144 67 148 71
rect 169 67 173 71
rect -41 55 -31 59
rect -41 33 -37 55
rect -41 29 -24 33
rect -41 -1 -37 29
rect -17 -1 -13 59
rect -1 53 3 59
rect -1 -1 3 48
rect 16 24 20 59
rect 16 20 24 24
rect 16 3 20 20
rect 40 18 44 59
rect 40 14 57 18
rect 27 6 33 10
rect 40 3 44 14
rect 64 6 68 59
rect 80 55 90 59
rect 104 55 114 59
rect 128 55 138 59
rect 152 55 162 59
rect 177 55 187 59
rect 80 32 84 55
rect 80 28 88 32
rect 16 -1 26 3
rect 40 -1 50 3
rect 64 2 73 6
rect 64 -1 68 2
rect 80 -1 84 28
rect 104 16 108 55
rect 104 12 121 16
rect 128 12 132 55
rect 152 51 156 55
rect 152 47 170 51
rect 104 -1 108 12
rect 128 8 145 12
rect 128 -1 132 8
rect 152 -1 156 47
rect 177 24 181 55
rect 177 20 191 24
rect 177 -1 181 20
rect -49 -9 -45 -5
rect -33 -9 -29 -5
rect -25 -9 -21 -5
rect -9 -9 -5 -5
rect 8 -9 12 -5
rect 32 -9 36 -5
rect 56 -9 60 -5
rect 72 -9 76 -5
rect 88 -9 92 -5
rect 96 -9 100 -5
rect 112 -9 116 -5
rect 120 -9 124 -5
rect 136 -9 140 -5
rect 144 -9 148 -5
rect 160 -9 164 -5
rect 169 -9 173 -5
rect 185 -9 189 -5
rect -49 -10 189 -9
rect -45 -14 -41 -10
rect -37 -14 -33 -10
rect -29 -12 72 -10
rect -29 -14 -25 -12
rect -49 -16 -25 -14
rect -21 -16 -17 -12
rect -13 -16 -9 -12
rect -5 -16 -1 -12
rect 3 -16 8 -12
rect 12 -16 19 -12
rect 23 -16 32 -12
rect 36 -16 43 -12
rect 47 -16 56 -12
rect 60 -16 64 -12
rect 68 -14 72 -12
rect 76 -14 80 -10
rect 84 -14 88 -10
rect 92 -14 96 -10
rect 100 -14 104 -10
rect 108 -14 112 -10
rect 116 -14 120 -10
rect 124 -14 128 -10
rect 132 -14 136 -10
rect 140 -14 144 -10
rect 148 -14 152 -10
rect 156 -14 160 -10
rect 164 -14 169 -10
rect 173 -14 177 -10
rect 181 -14 185 -10
rect 68 -16 189 -14
rect -49 -17 189 -16
<< m2contact >>
rect -1 48 4 53
rect -13 39 -8 44
rect 24 20 29 25
rect 88 28 93 33
<< pm12contact >>
rect 8 48 13 53
rect 47 6 52 11
rect 87 47 92 52
rect 135 20 140 25
rect 96 6 101 11
rect 159 28 164 33
rect 184 39 189 44
<< metal2 >>
rect 4 48 8 52
rect 13 48 87 52
rect -8 39 184 43
rect 93 29 159 33
rect 29 20 135 24
rect 52 6 96 10
<< labels >>
rlabel polycontact -48 48 -44 52 1 S2
rlabel polycontact -34 48 -30 52 1 RST
rlabel polycontact -8 49 -4 53 1 S1
rlabel metal1 23 6 37 10 1 T
rlabel pm12contact 47 6 52 11 1 S0
rlabel polycontact 111 7 115 8 1 REQ
rlabel metal1 187 20 191 24 7 N1
rlabel metal1 -28 71 -28 79 1 VDD
rlabel metal1 -28 -17 -28 -9 1 GND
<< end >>
