magic
tech scmos
timestamp 1732217075
<< nwell >>
rect -5 73 292 101
<< ntransistor >>
rect 7 15 9 19
rect 13 15 15 19
rect 31 15 33 19
rect 47 15 49 19
rect 55 15 57 19
rect 71 15 73 19
rect 79 15 81 19
rect 95 15 97 19
rect 101 15 103 19
rect 119 15 121 19
rect 135 15 137 19
rect 143 15 145 19
rect 159 15 161 19
rect 167 15 169 19
rect 183 15 185 19
rect 189 15 191 19
rect 207 15 209 19
rect 223 15 225 19
rect 231 15 233 19
rect 247 15 249 19
rect 255 15 257 19
rect 273 15 275 19
rect 279 15 281 19
<< ptransistor >>
rect 7 79 9 87
rect 15 79 17 87
rect 31 79 33 87
rect 49 79 51 87
rect 55 79 57 87
rect 73 79 75 87
rect 79 79 81 87
rect 95 79 97 87
rect 103 79 105 87
rect 119 79 121 87
rect 137 79 139 87
rect 143 79 145 87
rect 161 79 163 87
rect 167 79 169 87
rect 183 79 185 87
rect 191 79 193 87
rect 207 79 209 87
rect 225 79 227 87
rect 231 79 233 87
rect 249 79 251 87
rect 255 79 257 87
rect 271 79 273 87
rect 279 79 281 87
<< ndiffusion >>
rect 6 15 7 19
rect 9 15 13 19
rect 15 15 16 19
rect 30 15 31 19
rect 33 15 34 19
rect 46 15 47 19
rect 49 15 50 19
rect 54 15 55 19
rect 57 15 58 19
rect 70 15 71 19
rect 73 15 74 19
rect 78 15 79 19
rect 81 15 82 19
rect 94 15 95 19
rect 97 15 101 19
rect 103 15 104 19
rect 118 15 119 19
rect 121 15 122 19
rect 134 15 135 19
rect 137 15 138 19
rect 142 15 143 19
rect 145 15 146 19
rect 158 15 159 19
rect 161 15 162 19
rect 166 15 167 19
rect 169 15 170 19
rect 182 15 183 19
rect 185 15 189 19
rect 191 15 192 19
rect 206 15 207 19
rect 209 15 210 19
rect 222 15 223 19
rect 225 15 226 19
rect 230 15 231 19
rect 233 15 234 19
rect 246 15 247 19
rect 249 15 250 19
rect 254 15 255 19
rect 257 15 258 19
rect 272 15 273 19
rect 275 15 279 19
rect 281 15 282 19
<< pdiffusion >>
rect 6 79 7 87
rect 9 79 10 87
rect 14 79 15 87
rect 17 79 18 87
rect 30 79 31 87
rect 33 79 34 87
rect 48 79 49 87
rect 51 79 55 87
rect 57 79 58 87
rect 72 79 73 87
rect 75 79 79 87
rect 81 79 82 87
rect 94 79 95 87
rect 97 79 98 87
rect 102 79 103 87
rect 105 79 106 87
rect 118 79 119 87
rect 121 79 122 87
rect 136 79 137 87
rect 139 79 143 87
rect 145 79 146 87
rect 160 79 161 87
rect 163 79 167 87
rect 169 79 170 87
rect 182 79 183 87
rect 185 79 186 87
rect 190 79 191 87
rect 193 79 194 87
rect 206 79 207 87
rect 209 79 210 87
rect 224 79 225 87
rect 227 79 231 87
rect 233 79 234 87
rect 248 79 249 87
rect 251 79 255 87
rect 257 79 258 87
rect 270 79 271 87
rect 273 79 274 87
rect 278 79 279 87
rect 281 79 282 87
<< ndcontact >>
rect 2 15 6 19
rect 16 15 20 19
rect 26 15 30 19
rect 34 15 38 19
rect 42 15 46 19
rect 50 15 54 19
rect 58 15 62 19
rect 66 15 70 19
rect 74 15 78 19
rect 82 15 86 19
rect 90 15 94 19
rect 104 15 108 19
rect 114 15 118 19
rect 122 15 126 19
rect 130 15 134 19
rect 138 15 142 19
rect 146 15 150 19
rect 154 15 158 19
rect 162 15 166 19
rect 170 15 174 19
rect 178 15 182 19
rect 192 15 196 19
rect 202 15 206 19
rect 210 15 214 19
rect 218 15 222 19
rect 226 15 230 19
rect 234 15 238 19
rect 242 15 246 19
rect 250 15 254 19
rect 258 15 262 19
rect 268 15 272 19
rect 282 15 286 19
<< pdcontact >>
rect 2 79 6 87
rect 10 79 14 87
rect 18 79 22 87
rect 26 79 30 87
rect 34 79 38 87
rect 44 79 48 87
rect 58 79 62 87
rect 68 79 72 87
rect 82 79 86 87
rect 90 79 94 87
rect 98 79 102 87
rect 106 79 110 87
rect 114 79 118 87
rect 122 79 126 87
rect 132 79 136 87
rect 146 79 150 87
rect 156 79 160 87
rect 170 79 174 87
rect 178 79 182 87
rect 186 79 190 87
rect 194 79 198 87
rect 202 79 206 87
rect 210 79 214 87
rect 220 79 224 87
rect 234 79 238 87
rect 244 79 248 87
rect 258 79 262 87
rect 266 79 270 87
rect 274 79 278 87
rect 282 79 286 87
<< psubstratepcontact >>
rect 2 4 6 8
rect 13 4 17 8
rect 26 4 30 8
rect 34 4 38 8
rect 42 4 46 8
rect 50 4 54 8
rect 58 4 62 8
rect 66 4 70 8
rect 74 4 78 8
rect 82 4 86 8
rect 90 4 94 8
rect 101 4 105 8
rect 114 4 118 8
rect 122 4 126 8
rect 130 4 134 8
rect 138 4 142 8
rect 146 4 150 8
rect 154 4 158 8
rect 162 4 166 8
rect 170 4 174 8
rect 178 4 182 8
rect 189 4 193 8
rect 202 4 206 8
rect 210 4 214 8
rect 218 4 222 8
rect 226 4 230 8
rect 234 4 238 8
rect 242 4 246 8
rect 250 4 254 8
rect 258 4 262 8
rect 271 4 275 8
rect 282 4 286 8
<< nsubstratencontact >>
rect 2 94 6 98
rect 10 94 14 98
rect 18 94 22 98
rect 26 94 30 98
rect 34 94 38 98
rect 44 94 48 98
rect 58 94 62 98
rect 68 94 72 98
rect 82 94 86 98
rect 90 94 94 98
rect 98 94 102 98
rect 106 94 110 98
rect 114 94 118 98
rect 122 94 126 98
rect 132 94 136 98
rect 146 94 150 98
rect 156 94 160 98
rect 170 94 174 98
rect 178 94 182 98
rect 186 94 190 98
rect 194 94 198 98
rect 202 94 206 98
rect 210 94 214 98
rect 220 94 224 98
rect 234 94 238 98
rect 244 94 248 98
rect 258 94 262 98
rect 266 94 270 98
rect 274 94 278 98
rect 282 94 286 98
<< polysilicon >>
rect 7 87 9 90
rect 15 87 17 90
rect 31 87 33 90
rect 49 87 51 90
rect 55 87 57 90
rect 73 87 75 90
rect 79 87 81 90
rect 95 87 97 90
rect 103 87 105 90
rect 119 87 121 90
rect 137 87 139 90
rect 143 87 145 90
rect 161 87 163 90
rect 167 87 169 90
rect 183 87 185 90
rect 191 87 193 90
rect 207 87 209 90
rect 225 87 227 90
rect 231 87 233 90
rect 249 87 251 90
rect 255 87 257 90
rect 271 87 273 90
rect 279 87 281 90
rect 7 19 9 79
rect 15 27 17 79
rect 31 53 33 79
rect 49 54 51 79
rect 30 49 33 53
rect 13 25 17 27
rect 13 19 15 25
rect 31 19 33 49
rect 47 52 51 54
rect 47 19 49 52
rect 55 19 57 79
rect 73 48 75 79
rect 71 46 75 48
rect 71 19 73 46
rect 79 19 81 79
rect 95 19 97 79
rect 103 27 105 79
rect 119 41 121 79
rect 137 51 139 79
rect 135 49 139 51
rect 118 37 121 41
rect 101 25 105 27
rect 101 19 103 25
rect 119 19 121 37
rect 135 19 137 49
rect 143 19 145 79
rect 161 42 163 79
rect 159 40 163 42
rect 159 19 161 40
rect 167 19 169 79
rect 183 19 185 79
rect 191 27 193 79
rect 207 42 209 79
rect 225 50 227 79
rect 206 38 209 42
rect 189 25 193 27
rect 189 19 191 25
rect 207 19 209 38
rect 223 48 227 50
rect 223 19 225 48
rect 231 19 233 79
rect 249 44 251 79
rect 247 42 251 44
rect 247 19 249 42
rect 255 19 257 79
rect 271 26 273 79
rect 271 24 275 26
rect 273 19 275 24
rect 279 19 281 79
rect 7 12 9 15
rect 13 12 15 15
rect 31 12 33 15
rect 47 12 49 15
rect 55 12 57 15
rect 71 12 73 15
rect 79 12 81 15
rect 95 12 97 15
rect 101 12 103 15
rect 119 12 121 15
rect 135 12 137 15
rect 143 12 145 15
rect 159 12 161 15
rect 167 12 169 15
rect 183 12 185 15
rect 189 12 191 15
rect 207 12 209 15
rect 223 12 225 15
rect 231 12 233 15
rect 247 12 249 15
rect 255 12 257 15
rect 273 12 275 15
rect 279 12 281 15
<< polycontact >>
rect 26 49 30 53
rect 43 30 47 34
rect 57 30 61 34
rect 114 37 118 41
rect 131 30 135 34
rect 145 30 149 34
rect 202 38 206 42
rect 219 30 223 34
rect 233 30 237 34
<< metal1 >>
rect 2 98 286 99
rect 6 94 10 98
rect 14 94 18 98
rect 22 94 26 98
rect 30 94 34 98
rect 38 94 44 98
rect 48 94 58 98
rect 62 94 68 98
rect 72 94 82 98
rect 86 94 90 98
rect 94 94 98 98
rect 102 94 106 98
rect 110 94 114 98
rect 118 94 122 98
rect 126 94 132 98
rect 136 94 146 98
rect 150 94 156 98
rect 160 94 170 98
rect 174 94 178 98
rect 182 94 186 98
rect 190 94 194 98
rect 198 94 202 98
rect 206 94 210 98
rect 214 94 220 98
rect 224 94 234 98
rect 238 94 244 98
rect 248 94 258 98
rect 262 94 266 98
rect 270 94 274 98
rect 278 94 282 98
rect 2 91 286 94
rect 2 87 6 91
rect 18 87 22 91
rect 26 87 30 91
rect 58 87 62 91
rect 82 87 86 91
rect 10 34 14 79
rect 34 64 38 79
rect 90 87 94 91
rect 106 87 110 91
rect 114 87 118 91
rect 146 87 150 91
rect 170 87 174 91
rect 44 59 48 79
rect 26 34 30 49
rect 10 30 30 34
rect 34 34 38 59
rect 42 55 48 59
rect 68 57 72 79
rect 42 48 46 55
rect 66 53 72 57
rect 41 44 54 48
rect 41 43 46 44
rect 34 30 43 34
rect 10 29 22 30
rect 18 24 22 29
rect 16 21 22 24
rect 16 19 20 21
rect 34 19 38 30
rect 50 19 54 44
rect 66 34 70 53
rect 98 36 102 79
rect 114 36 118 37
rect 61 30 78 34
rect 98 31 106 36
rect 111 31 118 36
rect 122 34 126 79
rect 178 87 182 91
rect 194 87 198 91
rect 202 87 206 91
rect 234 87 238 91
rect 258 87 262 91
rect 132 56 136 79
rect 130 52 136 56
rect 130 42 134 52
rect 156 48 160 79
rect 154 44 160 48
rect 134 38 142 42
rect 74 19 78 30
rect 106 24 110 31
rect 104 21 110 24
rect 122 30 131 34
rect 104 19 108 21
rect 122 19 126 30
rect 138 19 142 38
rect 154 34 158 44
rect 186 36 190 79
rect 202 36 206 38
rect 149 30 166 34
rect 186 31 194 36
rect 199 32 206 36
rect 210 34 214 79
rect 266 87 270 91
rect 282 87 286 91
rect 220 56 224 79
rect 218 52 224 56
rect 244 54 248 79
rect 218 42 222 52
rect 242 49 248 54
rect 217 38 230 42
rect 217 37 222 38
rect 162 19 166 30
rect 194 24 198 31
rect 192 21 198 24
rect 210 30 219 34
rect 192 19 196 21
rect 210 19 214 30
rect 226 19 230 38
rect 242 34 246 49
rect 274 35 278 79
rect 237 30 254 34
rect 266 32 278 35
rect 250 19 254 30
rect 261 31 278 32
rect 261 27 270 31
rect 266 23 270 27
rect 266 21 272 23
rect 267 20 272 21
rect 268 19 272 20
rect 2 11 6 15
rect 26 11 30 15
rect 42 11 46 15
rect 58 11 62 15
rect 66 11 70 15
rect 82 11 86 15
rect 90 11 94 15
rect 114 11 118 15
rect 130 11 134 15
rect 146 11 150 15
rect 154 11 158 15
rect 170 11 174 15
rect 178 11 182 15
rect 202 11 206 15
rect 218 11 222 15
rect 234 11 238 15
rect 242 11 246 15
rect 258 11 262 15
rect 282 11 286 15
rect 2 8 286 11
rect 6 4 13 8
rect 17 4 26 8
rect 30 4 34 8
rect 38 4 42 8
rect 46 4 50 8
rect 54 4 58 8
rect 62 4 66 8
rect 70 4 74 8
rect 78 4 82 8
rect 86 4 90 8
rect 94 4 101 8
rect 105 4 114 8
rect 118 4 122 8
rect 126 4 130 8
rect 134 4 138 8
rect 142 4 146 8
rect 150 4 154 8
rect 158 4 162 8
rect 166 4 170 8
rect 174 4 178 8
rect 182 4 189 8
rect 193 4 202 8
rect 206 4 210 8
rect 214 4 218 8
rect 222 4 226 8
rect 230 4 234 8
rect 238 4 242 8
rect 246 4 250 8
rect 254 4 258 8
rect 262 4 271 8
rect 275 4 282 8
rect 2 3 286 4
<< m2contact >>
rect 34 59 39 64
rect 106 31 111 36
rect 194 31 199 36
<< pm12contact >>
rect 17 68 22 73
rect 81 68 86 73
rect 2 22 7 27
rect 105 68 110 73
rect 169 68 174 73
rect 66 22 71 27
rect 90 22 95 27
rect 193 68 198 73
rect 257 68 262 73
rect 266 51 271 56
rect 154 22 159 27
rect 178 22 183 27
rect 281 43 286 48
rect 242 22 247 27
<< ndm12contact >>
rect 129 37 134 42
<< metal2 >>
rect 22 68 81 73
rect 110 68 169 73
rect 198 68 257 73
rect 194 63 198 68
rect 39 59 198 63
rect 106 51 266 55
rect 106 36 110 51
rect 194 43 281 47
rect 134 37 176 42
rect 172 27 176 37
rect 194 36 198 43
rect 7 22 66 27
rect 95 22 154 27
rect 172 22 178 27
rect 183 22 242 27
<< labels >>
rlabel nwell 2 91 22 99 1 VDD
rlabel metal1 9 6 9 6 1 GND
rlabel metal1 44 45 44 47 1 Sum1
rlabel metal1 264 29 264 29 1 Cout
rlabel metal1 220 39 220 41 1 Sum2
rlabel pm12contact 2 23 2 27 1 A0
rlabel metal2 22 69 22 73 1 B0
rlabel metal2 110 69 110 73 1 B1
rlabel pm12contact 90 23 90 27 1 A1
<< end >>
