magic
tech scmos
timestamp 1732203366
<< nwell >>
rect -16 19 14 47
<< ntransistor >>
rect -5 -39 -3 -35
rect 3 -39 5 -35
<< ptransistor >>
rect -5 25 -3 33
rect 1 25 3 33
<< ndiffusion >>
rect -6 -39 -5 -35
rect -3 -39 -2 -35
rect 2 -39 3 -35
rect 5 -39 6 -35
<< pdiffusion >>
rect -6 25 -5 33
rect -3 25 1 33
rect 3 25 4 33
<< ndcontact >>
rect -10 -39 -6 -35
rect -2 -39 2 -35
rect 6 -39 10 -35
<< pdcontact >>
rect -10 25 -6 33
rect 4 25 8 33
<< psubstratepcontact >>
rect -10 -50 -6 -46
rect -2 -50 2 -46
rect 6 -51 10 -47
<< nsubstratencontact >>
rect -10 40 -6 44
rect 4 40 8 44
<< polysilicon >>
rect -5 33 -3 36
rect 1 33 3 36
rect -5 -35 -3 25
rect 1 -6 3 25
rect 1 -8 5 -6
rect 3 -35 5 -8
rect -5 -42 -3 -39
rect 3 -42 5 -39
<< polycontact >>
rect -9 -3 -5 1
rect 5 -27 9 -23
<< metal1 >>
rect -10 44 8 45
rect -6 40 4 44
rect -10 37 8 40
rect -10 33 -6 37
rect 4 3 8 25
rect 4 -1 10 3
rect 6 -4 10 -1
rect 6 -8 14 -4
rect 6 -12 10 -8
rect -2 -16 10 -12
rect -2 -35 2 -16
rect -10 -43 -6 -39
rect 6 -43 10 -39
rect -10 -46 10 -43
rect -6 -50 -2 -46
rect 2 -47 10 -46
rect 2 -50 6 -47
rect -10 -51 6 -50
<< labels >>
rlabel polycontact -9 -3 -5 1 1 A
rlabel polycontact 5 -27 9 -23 1 B
rlabel metal1 10 -8 14 -4 7 Y
rlabel metal1 -10 -51 10 -43 1 GND
rlabel nwell -10 37 8 45 1 VDD
<< end >>
