module sett_less_than(
	output [31:0] set_less_than,
	input less_than

);


	and and_0(set_less_than[0],less_than,1);
	and and_1(set_less_than[1],0 ,less_than);
	and and_2(set_less_than[2],0 ,less_than);
	and and_3(set_less_than[3],0 ,less_than);
	and and_4(set_less_than[4],0 ,less_than);
	and and_5(set_less_than[5],0 ,less_than);
	and and_6(set_less_than[6],0 ,less_than);
	and and_7(set_less_than[7],0 ,less_than);
	and and_8(set_less_than[8],0 ,less_than);
	and and_9(set_less_than[9],0 ,less_than);
	and and_10(set_less_than[10],0 ,less_than);
	and and_11(set_less_than[11],0 ,less_than);
	and and_12(set_less_than[12],0 ,less_than);
	and and_13(set_less_than[13],0 ,less_than);
	and and_14(set_less_than[14],0 ,less_than);
	and and_15(set_less_than[15],0 ,less_than);
	and and_16(set_less_than[16],0 ,less_than);
	and and_17(set_less_than[17],0 ,less_than);
	and and_18(set_less_than[18],0 ,less_than);
	and and_19(set_less_than[19],0 ,less_than);
	and and_20(set_less_than[20],0 ,less_than);
	and and_21(set_less_than[21],0 ,less_than);
	and and_22(set_less_than[22],0 ,less_than);
	and and_23(set_less_than[23],0 ,less_than);
	and and_24(set_less_than[24],0 ,less_than);
	and and_25(set_less_than[25],0 ,less_than);
	and and_26(set_less_than[26],0 ,less_than);
	and and_27(set_less_than[27],0 ,less_than);
	and and_28(set_less_than[28],0 ,less_than);
	and and_29(set_less_than[29],0 ,less_than);
	and and_30(set_less_than[30],0 ,less_than);
	and and_31(set_less_than[31],0 ,less_than);


	

endmodule 