module generator_4bit(
	
	
	
	input in_0[3:0];
	input in_1[3:0];
);








endmodule 