magic
tech scmos
timestamp 1736883192
<< nwell >>
rect -181 65 482 93
rect 56 -75 77 -74
rect -191 -107 593 -75
<< ntransistor >>
rect -172 7 -170 11
rect -164 7 -162 11
rect -140 7 -138 11
rect -117 7 -115 11
rect -94 7 -92 11
rect -86 7 -84 11
rect -70 7 -68 11
rect -62 7 -60 11
rect -6 7 -4 11
rect 2 7 4 11
rect 18 7 20 11
rect 34 7 36 11
rect 51 7 53 11
rect 57 7 59 11
rect 89 7 91 11
rect 113 7 115 11
rect 119 7 121 11
rect 137 7 139 11
rect 153 7 155 11
rect 161 7 163 11
rect 177 7 179 11
rect 185 7 187 11
rect 201 7 203 11
rect 209 7 211 11
rect 225 7 227 11
rect 233 7 235 11
rect 250 7 252 11
rect 258 7 260 11
rect 290 7 292 11
rect 296 7 298 11
rect 326 7 328 11
rect 332 7 334 11
rect 350 7 352 11
rect 366 7 368 11
rect 374 7 376 11
rect 390 7 392 11
rect 398 7 400 11
rect 414 7 416 11
rect 422 7 424 11
rect 438 7 440 11
rect 446 7 448 11
rect 463 7 465 11
rect 471 7 473 11
rect -180 -12 -178 -8
rect -158 -14 -156 -10
rect -132 -12 -130 -8
rect -126 -12 -124 -8
rect -118 -12 -116 -8
rect -88 -12 -86 -8
rect -80 -12 -78 -8
rect -74 -12 -72 -8
rect -56 -12 -54 -8
rect -32 -14 -30 -10
rect -10 -12 -8 -8
rect -4 -12 -2 -8
rect 4 -12 6 -8
rect 34 -12 36 -8
rect 42 -12 44 -8
rect 48 -12 50 -8
rect 82 -12 84 -8
rect 88 -12 90 -8
rect 96 -12 98 -8
rect 128 -12 130 -8
rect 136 -12 138 -8
rect 142 -12 144 -8
rect 164 -14 166 -10
rect 188 -12 190 -8
rect 206 -12 208 -8
rect 212 -12 214 -8
rect 220 -12 222 -8
rect 250 -12 252 -8
rect 258 -12 260 -8
rect 264 -12 266 -8
rect 290 -14 292 -10
rect 312 -12 314 -8
rect 349 -12 351 -8
rect 355 -12 357 -8
rect 363 -12 365 -8
rect 393 -12 395 -8
rect 401 -12 403 -8
rect 407 -12 409 -8
rect 429 -14 431 -10
rect 453 -12 455 -8
rect 471 -12 473 -8
rect 477 -12 479 -8
rect 485 -12 487 -8
rect 515 -12 517 -8
rect 523 -12 525 -8
rect 529 -12 531 -8
rect 558 -14 560 -10
rect 580 -12 582 -8
<< ptransistor >>
rect -170 71 -168 79
rect -164 71 -162 79
rect -140 71 -138 79
rect -117 71 -115 79
rect -94 71 -92 79
rect -88 71 -86 79
rect -68 71 -66 79
rect -62 71 -60 79
rect -6 71 -4 79
rect 0 71 2 79
rect 18 71 20 79
rect 34 71 36 79
rect 51 71 53 79
rect 59 71 61 79
rect 89 71 91 79
rect 113 71 115 79
rect 121 71 123 79
rect 137 71 139 79
rect 153 71 155 79
rect 159 71 161 79
rect 177 71 179 79
rect 183 71 185 79
rect 201 71 203 79
rect 207 71 209 79
rect 225 71 227 79
rect 231 71 233 79
rect 250 71 252 79
rect 256 71 258 79
rect 290 71 292 79
rect 298 71 300 79
rect 326 71 328 79
rect 334 71 336 79
rect 350 71 352 79
rect 366 71 368 79
rect 372 71 374 79
rect 390 71 392 79
rect 396 71 398 79
rect 414 71 416 79
rect 420 71 422 79
rect 438 71 440 79
rect 444 71 446 79
rect 463 71 465 79
rect 469 71 471 79
rect -180 -89 -178 -81
rect -158 -89 -156 -81
rect -132 -89 -130 -81
rect -124 -89 -122 -81
rect -116 -89 -114 -81
rect -90 -89 -88 -81
rect -82 -89 -80 -81
rect -74 -89 -72 -81
rect -56 -89 -54 -81
rect -32 -89 -30 -81
rect -10 -89 -8 -81
rect -2 -89 0 -81
rect 6 -89 8 -81
rect 32 -89 34 -81
rect 40 -89 42 -81
rect 48 -89 50 -81
rect 82 -89 84 -81
rect 90 -89 92 -81
rect 98 -89 100 -81
rect 126 -89 128 -81
rect 134 -89 136 -81
rect 142 -89 144 -81
rect 164 -89 166 -81
rect 188 -89 190 -81
rect 206 -89 208 -81
rect 214 -89 216 -81
rect 222 -89 224 -81
rect 248 -89 250 -81
rect 256 -89 258 -81
rect 264 -89 266 -81
rect 290 -89 292 -81
rect 312 -89 314 -81
rect 349 -89 351 -81
rect 357 -89 359 -81
rect 365 -89 367 -81
rect 391 -89 393 -81
rect 399 -89 401 -81
rect 407 -89 409 -81
rect 429 -89 431 -81
rect 453 -89 455 -81
rect 471 -89 473 -81
rect 479 -89 481 -81
rect 487 -89 489 -81
rect 513 -89 515 -81
rect 521 -89 523 -81
rect 529 -89 531 -81
rect 558 -89 560 -81
rect 580 -89 582 -81
<< ndiffusion >>
rect -173 7 -172 11
rect -170 7 -169 11
rect -165 7 -164 11
rect -162 7 -161 11
rect -141 7 -140 11
rect -138 7 -137 11
rect -118 7 -117 11
rect -115 7 -114 11
rect -95 7 -94 11
rect -92 7 -91 11
rect -87 7 -86 11
rect -84 7 -83 11
rect -71 7 -70 11
rect -68 7 -67 11
rect -63 7 -62 11
rect -60 7 -59 11
rect -7 7 -6 11
rect -4 7 -3 11
rect 1 7 2 11
rect 4 7 5 11
rect 17 7 18 11
rect 20 7 21 11
rect 33 7 34 11
rect 36 7 37 11
rect 50 7 51 11
rect 53 7 57 11
rect 59 7 60 11
rect 88 7 89 11
rect 91 7 92 11
rect 112 7 113 11
rect 115 7 119 11
rect 121 7 122 11
rect 136 7 137 11
rect 139 7 140 11
rect 152 7 153 11
rect 155 7 156 11
rect 160 7 161 11
rect 163 7 164 11
rect 176 7 177 11
rect 179 7 180 11
rect 184 7 185 11
rect 187 7 188 11
rect 200 7 201 11
rect 203 7 204 11
rect 208 7 209 11
rect 211 7 212 11
rect 224 7 225 11
rect 227 7 228 11
rect 232 7 233 11
rect 235 7 236 11
rect 249 7 250 11
rect 252 7 253 11
rect 257 7 258 11
rect 260 7 261 11
rect 289 7 290 11
rect 292 7 296 11
rect 298 7 299 11
rect 325 7 326 11
rect 328 7 332 11
rect 334 7 335 11
rect 349 7 350 11
rect 352 7 353 11
rect 365 7 366 11
rect 368 7 369 11
rect 373 7 374 11
rect 376 7 377 11
rect 389 7 390 11
rect 392 7 393 11
rect 397 7 398 11
rect 400 7 401 11
rect 413 7 414 11
rect 416 7 417 11
rect 421 7 422 11
rect 424 7 425 11
rect 437 7 438 11
rect 440 7 441 11
rect 445 7 446 11
rect 448 7 449 11
rect 462 7 463 11
rect 465 7 466 11
rect 470 7 471 11
rect 473 7 474 11
rect -181 -12 -180 -8
rect -178 -12 -177 -8
rect -159 -14 -158 -10
rect -156 -14 -155 -10
rect -133 -12 -132 -8
rect -130 -12 -126 -8
rect -124 -12 -123 -8
rect -119 -12 -118 -8
rect -116 -12 -115 -8
rect -89 -12 -88 -8
rect -86 -12 -85 -8
rect -81 -12 -80 -8
rect -78 -12 -74 -8
rect -72 -12 -71 -8
rect -57 -12 -56 -8
rect -54 -12 -53 -8
rect -33 -14 -32 -10
rect -30 -14 -29 -10
rect -11 -12 -10 -8
rect -8 -12 -4 -8
rect -2 -12 -1 -8
rect 3 -12 4 -8
rect 6 -12 7 -8
rect 33 -12 34 -8
rect 36 -12 37 -8
rect 41 -12 42 -8
rect 44 -12 48 -8
rect 50 -12 51 -8
rect 81 -12 82 -8
rect 84 -12 88 -8
rect 90 -12 91 -8
rect 95 -12 96 -8
rect 98 -12 99 -8
rect 127 -12 128 -8
rect 130 -12 131 -8
rect 135 -12 136 -8
rect 138 -12 142 -8
rect 144 -12 145 -8
rect 163 -14 164 -10
rect 166 -14 167 -10
rect 187 -12 188 -8
rect 190 -12 191 -8
rect 205 -12 206 -8
rect 208 -12 212 -8
rect 214 -12 215 -8
rect 219 -12 220 -8
rect 222 -12 223 -8
rect 249 -12 250 -8
rect 252 -12 253 -8
rect 257 -12 258 -8
rect 260 -12 264 -8
rect 266 -12 267 -8
rect 289 -14 290 -10
rect 292 -14 293 -10
rect 311 -12 312 -8
rect 314 -12 315 -8
rect 348 -12 349 -8
rect 351 -12 355 -8
rect 357 -12 358 -8
rect 362 -12 363 -8
rect 365 -12 366 -8
rect 392 -12 393 -8
rect 395 -12 396 -8
rect 400 -12 401 -8
rect 403 -12 407 -8
rect 409 -12 410 -8
rect 428 -14 429 -10
rect 431 -14 432 -10
rect 452 -12 453 -8
rect 455 -12 456 -8
rect 470 -12 471 -8
rect 473 -12 477 -8
rect 479 -12 480 -8
rect 484 -12 485 -8
rect 487 -12 488 -8
rect 514 -12 515 -8
rect 517 -12 518 -8
rect 522 -12 523 -8
rect 525 -12 529 -8
rect 531 -12 532 -8
rect 557 -14 558 -10
rect 560 -14 561 -10
rect 579 -12 580 -8
rect 582 -12 583 -8
<< pdiffusion >>
rect -171 71 -170 79
rect -168 71 -164 79
rect -162 71 -161 79
rect -141 71 -140 79
rect -138 71 -137 79
rect -118 71 -117 79
rect -115 71 -114 79
rect -95 71 -94 79
rect -92 71 -88 79
rect -86 71 -85 79
rect -69 71 -68 79
rect -66 71 -62 79
rect -60 71 -59 79
rect -7 71 -6 79
rect -4 71 0 79
rect 2 71 3 79
rect 17 71 18 79
rect 20 71 21 79
rect 33 71 34 79
rect 36 71 37 79
rect 50 71 51 79
rect 53 71 54 79
rect 58 71 59 79
rect 61 71 62 79
rect 88 71 89 79
rect 91 71 92 79
rect 112 71 113 79
rect 115 71 116 79
rect 120 71 121 79
rect 123 71 124 79
rect 136 71 137 79
rect 139 71 140 79
rect 152 71 153 79
rect 155 71 159 79
rect 161 71 162 79
rect 176 71 177 79
rect 179 71 183 79
rect 185 71 186 79
rect 200 71 201 79
rect 203 71 207 79
rect 209 71 210 79
rect 224 71 225 79
rect 227 71 231 79
rect 233 71 234 79
rect 249 71 250 79
rect 252 71 256 79
rect 258 71 259 79
rect 289 71 290 79
rect 292 71 293 79
rect 297 71 298 79
rect 300 71 301 79
rect 325 71 326 79
rect 328 71 329 79
rect 333 71 334 79
rect 336 71 337 79
rect 349 71 350 79
rect 352 71 353 79
rect 365 71 366 79
rect 368 71 372 79
rect 374 71 375 79
rect 389 71 390 79
rect 392 71 396 79
rect 398 71 399 79
rect 413 71 414 79
rect 416 71 420 79
rect 422 71 423 79
rect 437 71 438 79
rect 440 71 444 79
rect 446 71 447 79
rect 462 71 463 79
rect 465 71 469 79
rect 471 71 472 79
rect -181 -89 -180 -81
rect -178 -89 -177 -81
rect -159 -89 -158 -81
rect -156 -89 -155 -81
rect -133 -89 -132 -81
rect -130 -89 -129 -81
rect -125 -89 -124 -81
rect -122 -89 -121 -81
rect -117 -89 -116 -81
rect -114 -89 -113 -81
rect -91 -89 -90 -81
rect -88 -89 -87 -81
rect -83 -89 -82 -81
rect -80 -89 -79 -81
rect -75 -89 -74 -81
rect -72 -89 -71 -81
rect -57 -89 -56 -81
rect -54 -89 -53 -81
rect -33 -89 -32 -81
rect -30 -89 -29 -81
rect -11 -89 -10 -81
rect -8 -89 -7 -81
rect -3 -89 -2 -81
rect 0 -89 1 -81
rect 5 -89 6 -81
rect 8 -89 9 -81
rect 31 -89 32 -81
rect 34 -89 35 -81
rect 39 -89 40 -81
rect 42 -89 43 -81
rect 47 -89 48 -81
rect 50 -89 51 -81
rect 81 -89 82 -81
rect 84 -89 85 -81
rect 89 -89 90 -81
rect 92 -89 93 -81
rect 97 -89 98 -81
rect 100 -89 101 -81
rect 125 -89 126 -81
rect 128 -89 129 -81
rect 133 -89 134 -81
rect 136 -89 137 -81
rect 141 -89 142 -81
rect 144 -89 145 -81
rect 163 -89 164 -81
rect 166 -89 167 -81
rect 187 -89 188 -81
rect 190 -89 191 -81
rect 205 -89 206 -81
rect 208 -89 209 -81
rect 213 -89 214 -81
rect 216 -89 217 -81
rect 221 -89 222 -81
rect 224 -89 225 -81
rect 247 -89 248 -81
rect 250 -89 251 -81
rect 255 -89 256 -81
rect 258 -89 259 -81
rect 263 -89 264 -81
rect 266 -89 267 -81
rect 289 -89 290 -81
rect 292 -89 293 -81
rect 311 -89 312 -81
rect 314 -89 315 -81
rect 348 -89 349 -81
rect 351 -89 352 -81
rect 356 -89 357 -81
rect 359 -89 360 -81
rect 364 -89 365 -81
rect 367 -89 368 -81
rect 390 -89 391 -81
rect 393 -89 394 -81
rect 398 -89 399 -81
rect 401 -89 402 -81
rect 406 -89 407 -81
rect 409 -89 410 -81
rect 428 -89 429 -81
rect 431 -89 432 -81
rect 452 -89 453 -81
rect 455 -89 456 -81
rect 470 -89 471 -81
rect 473 -89 474 -81
rect 478 -89 479 -81
rect 481 -89 482 -81
rect 486 -89 487 -81
rect 489 -89 490 -81
rect 512 -89 513 -81
rect 515 -89 516 -81
rect 520 -89 521 -81
rect 523 -89 524 -81
rect 528 -89 529 -81
rect 531 -89 532 -81
rect 557 -89 558 -81
rect 560 -89 561 -81
rect 579 -89 580 -81
rect 582 -89 583 -81
<< ndcontact >>
rect -177 7 -173 11
rect -169 7 -165 11
rect -161 7 -157 11
rect -145 7 -141 11
rect -137 7 -133 11
rect -122 7 -118 11
rect -114 7 -110 11
rect -99 7 -95 11
rect -91 7 -87 11
rect -83 7 -79 11
rect -75 7 -71 11
rect -67 7 -63 11
rect -59 7 -55 11
rect -11 7 -7 11
rect -3 7 1 11
rect 5 7 9 11
rect 13 7 17 11
rect 21 7 25 11
rect 29 7 33 11
rect 37 7 41 11
rect 46 7 50 11
rect 60 7 64 11
rect 84 7 88 11
rect 92 7 96 11
rect 108 7 112 11
rect 122 7 126 11
rect 132 7 136 11
rect 140 7 144 11
rect 148 7 152 11
rect 156 7 160 11
rect 164 7 168 11
rect 172 7 176 11
rect 180 7 184 11
rect 188 7 192 11
rect 196 7 200 11
rect 204 7 208 11
rect 212 7 216 11
rect 220 7 224 11
rect 228 7 232 11
rect 236 7 240 11
rect 245 7 249 11
rect 253 7 257 11
rect 261 7 265 11
rect 285 7 289 11
rect 299 7 303 11
rect 321 7 325 11
rect 335 7 339 11
rect 345 7 349 11
rect 353 7 357 11
rect 361 7 365 11
rect 369 7 373 11
rect 377 7 381 11
rect 385 7 389 11
rect 393 7 397 11
rect 401 7 405 11
rect 409 7 413 11
rect 417 7 421 11
rect 425 7 429 11
rect 433 7 437 11
rect 441 7 445 11
rect 449 7 453 11
rect 458 7 462 11
rect 466 7 470 11
rect 474 7 478 11
rect -185 -12 -181 -8
rect -177 -12 -173 -8
rect -163 -14 -159 -10
rect -155 -14 -151 -10
rect -137 -12 -133 -8
rect -123 -12 -119 -8
rect -115 -12 -111 -8
rect -93 -12 -89 -8
rect -85 -12 -81 -8
rect -71 -12 -67 -8
rect -61 -12 -57 -8
rect -53 -12 -49 -8
rect -37 -14 -33 -10
rect -29 -14 -25 -10
rect -15 -12 -11 -8
rect -1 -12 3 -8
rect 7 -12 11 -8
rect 29 -12 33 -8
rect 37 -12 41 -8
rect 51 -12 55 -8
rect 77 -12 81 -8
rect 91 -12 95 -8
rect 99 -12 103 -8
rect 123 -12 127 -8
rect 131 -12 135 -8
rect 145 -12 149 -8
rect 159 -14 163 -10
rect 167 -14 171 -10
rect 183 -12 187 -8
rect 191 -12 195 -8
rect 201 -12 205 -8
rect 215 -12 219 -8
rect 223 -12 227 -8
rect 245 -12 249 -8
rect 253 -12 257 -8
rect 267 -12 271 -8
rect 285 -14 289 -10
rect 293 -14 297 -10
rect 307 -12 311 -8
rect 315 -12 319 -8
rect 344 -12 348 -8
rect 358 -12 362 -8
rect 366 -12 370 -8
rect 388 -12 392 -8
rect 396 -12 400 -8
rect 410 -12 414 -8
rect 424 -14 428 -10
rect 432 -14 436 -10
rect 448 -12 452 -8
rect 456 -12 460 -8
rect 466 -12 470 -8
rect 480 -12 484 -8
rect 488 -12 492 -8
rect 510 -12 514 -8
rect 518 -12 522 -8
rect 532 -12 536 -8
rect 553 -14 557 -10
rect 561 -14 565 -10
rect 575 -12 579 -8
rect 583 -12 587 -8
<< pdcontact >>
rect -175 71 -171 79
rect -161 71 -157 79
rect -145 71 -141 79
rect -137 71 -133 79
rect -122 71 -118 79
rect -114 71 -110 79
rect -99 71 -95 79
rect -85 71 -81 79
rect -73 71 -69 79
rect -59 71 -55 79
rect -11 71 -7 79
rect 3 71 7 79
rect 13 71 17 79
rect 21 71 25 79
rect 29 71 33 79
rect 37 71 41 79
rect 46 71 50 79
rect 54 71 58 79
rect 62 71 66 79
rect 84 71 88 79
rect 92 71 96 79
rect 108 71 112 79
rect 116 71 120 79
rect 124 71 128 79
rect 132 71 136 79
rect 140 71 144 79
rect 148 71 152 79
rect 162 71 166 79
rect 172 71 176 79
rect 186 71 190 79
rect 196 71 200 79
rect 210 71 214 79
rect 220 71 224 79
rect 234 71 238 79
rect 245 71 249 79
rect 259 71 263 79
rect 285 71 289 79
rect 293 71 297 79
rect 301 71 305 79
rect 321 71 325 79
rect 329 71 333 79
rect 337 71 341 79
rect 345 71 349 79
rect 353 71 357 79
rect 361 71 365 79
rect 375 71 379 79
rect 385 71 389 79
rect 399 71 403 79
rect 409 71 413 79
rect 423 71 427 79
rect 433 71 437 79
rect 447 71 451 79
rect 458 71 462 79
rect 472 71 476 79
rect -185 -89 -181 -81
rect -177 -89 -173 -81
rect -163 -89 -159 -81
rect -155 -89 -151 -81
rect -137 -89 -133 -81
rect -129 -89 -125 -81
rect -121 -89 -117 -81
rect -113 -89 -109 -81
rect -95 -89 -91 -81
rect -87 -89 -83 -81
rect -79 -89 -75 -81
rect -71 -89 -67 -81
rect -61 -89 -57 -81
rect -53 -89 -49 -81
rect -37 -89 -33 -81
rect -29 -89 -25 -81
rect -15 -89 -11 -81
rect -7 -89 -3 -81
rect 1 -89 5 -81
rect 9 -89 13 -81
rect 27 -89 31 -81
rect 35 -89 39 -81
rect 43 -89 47 -81
rect 51 -89 55 -81
rect 77 -89 81 -81
rect 85 -89 89 -81
rect 93 -89 97 -81
rect 101 -89 105 -81
rect 121 -89 125 -81
rect 129 -89 133 -81
rect 137 -89 141 -81
rect 145 -89 149 -81
rect 159 -89 163 -81
rect 167 -89 171 -81
rect 183 -89 187 -81
rect 191 -89 195 -81
rect 201 -89 205 -81
rect 209 -89 213 -81
rect 217 -89 221 -81
rect 225 -89 229 -81
rect 243 -89 247 -81
rect 251 -89 255 -81
rect 259 -89 263 -81
rect 267 -89 271 -81
rect 285 -89 289 -81
rect 293 -89 297 -81
rect 307 -89 311 -81
rect 315 -89 319 -81
rect 344 -89 348 -81
rect 352 -89 356 -81
rect 360 -89 364 -81
rect 368 -89 372 -81
rect 386 -89 390 -81
rect 394 -89 398 -81
rect 402 -89 406 -81
rect 410 -89 414 -81
rect 424 -89 428 -81
rect 432 -89 436 -81
rect 448 -89 452 -81
rect 456 -89 460 -81
rect 466 -89 470 -81
rect 474 -89 478 -81
rect 482 -89 486 -81
rect 490 -89 494 -81
rect 508 -89 512 -81
rect 516 -89 520 -81
rect 524 -89 528 -81
rect 532 -89 536 -81
rect 553 -89 557 -81
rect 561 -89 565 -81
rect 575 -89 579 -81
rect 583 -89 587 -81
<< psubstratepdiff >>
rect -11 -4 -7 -2
rect 13 -4 17 -2
rect 21 -4 25 -2
rect 46 -4 50 -2
rect 57 -4 61 -2
rect 84 -4 88 -2
rect 108 -4 112 -2
rect 119 -4 123 -2
rect 134 -4 144 -2
rect 297 -4 300 -2
rect 321 -4 325 -2
rect 332 -4 336 -2
rect 353 -4 357 -2
<< psubstratepcontact >>
rect -185 -2 -181 2
rect -177 -2 -49 2
rect -37 -2 -33 2
rect -29 -2 -25 2
rect -15 -2 492 2
rect 510 -2 514 2
rect 518 -2 522 2
rect 532 -2 536 2
rect 553 -2 557 2
rect 561 -2 565 2
rect 575 -2 579 2
rect 583 -2 587 2
<< nsubstratencontact >>
rect -176 85 -172 89
rect -168 85 -164 89
rect -160 85 -156 89
rect -145 85 -141 89
rect -137 85 -133 89
rect -122 85 -118 89
rect -114 85 -110 89
rect -100 85 -96 89
rect -92 85 -88 89
rect -84 85 -80 89
rect -74 85 -70 89
rect -66 85 -62 89
rect -58 85 -54 89
rect -11 84 -7 88
rect 3 84 7 88
rect 13 86 17 90
rect 21 86 25 90
rect 29 86 33 90
rect 37 86 41 90
rect 46 86 50 90
rect 54 86 58 90
rect 62 86 66 90
rect 84 86 88 90
rect 92 86 96 90
rect 108 86 112 90
rect 116 86 120 90
rect 124 86 128 90
rect 132 86 136 90
rect 140 86 144 90
rect 148 84 152 88
rect 162 84 166 88
rect 172 84 176 88
rect 186 84 190 88
rect 196 84 200 88
rect 210 84 214 88
rect 220 84 224 88
rect 234 84 238 88
rect 245 84 249 88
rect 259 84 263 88
rect 285 86 289 90
rect 293 86 297 90
rect 301 86 305 90
rect 321 86 325 90
rect 329 86 333 90
rect 337 86 341 90
rect 345 86 349 90
rect 353 86 357 90
rect 361 84 365 88
rect 375 84 379 88
rect 385 84 389 88
rect 399 84 403 88
rect 409 84 413 88
rect 423 84 427 88
rect 433 84 437 88
rect 447 84 451 88
rect 458 84 462 88
rect 472 84 476 88
rect -185 -99 -181 -95
rect -177 -99 -173 -95
rect -163 -99 -159 -95
rect -155 -99 -151 -95
rect -137 -99 -133 -95
rect -129 -99 -125 -95
rect -121 -99 -117 -95
rect -113 -99 -109 -95
rect -95 -99 -91 -95
rect -87 -99 -83 -95
rect -79 -99 -75 -95
rect -71 -99 -67 -95
rect -37 -99 -33 -95
rect -29 -99 -25 -95
rect -15 -99 -11 -95
rect -7 -99 -3 -95
rect 1 -99 5 -95
rect 9 -99 13 -95
rect 27 -99 31 -95
rect 35 -99 39 -95
rect 43 -99 47 -95
rect 51 -99 55 -95
rect 77 -99 81 -95
rect 85 -99 89 -95
rect 93 -99 97 -95
rect 101 -99 105 -95
rect 121 -99 125 -95
rect 129 -99 133 -95
rect 137 -99 141 -95
rect 145 -99 149 -95
rect 159 -99 163 -95
rect 167 -99 171 -95
rect 201 -99 205 -95
rect 209 -99 213 -95
rect 217 -99 221 -95
rect 225 -99 229 -95
rect 243 -99 247 -95
rect 251 -99 255 -95
rect 259 -99 263 -95
rect 267 -99 271 -95
rect 285 -99 289 -95
rect 293 -99 297 -95
rect 307 -99 311 -95
rect 315 -99 319 -95
rect 344 -99 348 -95
rect 352 -99 356 -95
rect 360 -99 364 -95
rect 368 -99 372 -95
rect 386 -99 390 -95
rect 394 -99 398 -95
rect 402 -99 406 -95
rect 410 -99 414 -95
rect 424 -99 428 -95
rect 432 -99 436 -95
rect 466 -99 470 -95
rect 474 -99 478 -95
rect 482 -99 486 -95
rect 490 -99 494 -95
rect 508 -99 512 -95
rect 516 -99 520 -95
rect 524 -99 528 -95
rect 532 -99 536 -95
rect 553 -99 557 -95
rect 561 -99 565 -95
rect 575 -99 579 -95
rect 583 -99 587 -95
<< polysilicon >>
rect -170 79 -168 82
rect -164 79 -162 82
rect -140 79 -138 82
rect -117 79 -115 82
rect -94 79 -92 82
rect -88 79 -86 82
rect -68 79 -66 82
rect -62 79 -60 82
rect -6 79 -4 82
rect 0 79 2 82
rect 18 79 20 82
rect 34 79 36 82
rect 51 79 53 82
rect 59 79 61 82
rect 89 79 91 82
rect 113 79 115 82
rect 121 79 123 82
rect 137 79 139 82
rect 153 79 155 82
rect 159 79 161 82
rect 177 79 179 82
rect 183 79 185 82
rect 201 79 203 82
rect 207 79 209 82
rect 225 79 227 82
rect 231 79 233 82
rect 250 79 252 82
rect 256 79 258 82
rect 290 79 292 82
rect 298 79 300 82
rect 326 79 328 82
rect 334 79 336 82
rect 350 79 352 82
rect 366 79 368 82
rect 372 79 374 82
rect 390 79 392 82
rect 396 79 398 82
rect 414 79 416 82
rect 420 79 422 82
rect 438 79 440 82
rect 444 79 446 82
rect 463 79 465 82
rect 469 79 471 82
rect -170 52 -168 71
rect -172 50 -168 52
rect -172 11 -170 50
rect -164 11 -162 71
rect -140 11 -138 71
rect -117 11 -115 71
rect -94 11 -92 71
rect -88 58 -86 71
rect -68 68 -66 71
rect -70 66 -66 68
rect -88 56 -84 58
rect -86 11 -84 56
rect -70 11 -68 66
rect -62 11 -60 71
rect -6 11 -4 71
rect 0 70 2 71
rect 0 68 4 70
rect 2 11 4 68
rect 18 11 20 71
rect 34 11 36 71
rect 51 11 53 71
rect 59 15 61 71
rect 57 13 61 15
rect 57 11 59 13
rect 89 11 91 71
rect 113 11 115 71
rect 121 15 123 71
rect 119 13 123 15
rect 119 11 121 13
rect 137 11 139 71
rect 153 11 155 71
rect 159 70 161 71
rect 159 68 163 70
rect 161 11 163 68
rect 177 11 179 71
rect 183 70 185 71
rect 183 68 187 70
rect 185 11 187 68
rect 201 11 203 71
rect 207 70 209 71
rect 207 68 211 70
rect 209 11 211 68
rect 225 11 227 71
rect 231 70 233 71
rect 231 68 235 70
rect 233 11 235 68
rect 250 11 252 71
rect 256 70 258 71
rect 256 68 260 70
rect 258 11 260 68
rect 290 11 292 71
rect 298 15 300 71
rect 296 13 300 15
rect 296 11 298 13
rect 326 11 328 71
rect 334 15 336 71
rect 332 13 336 15
rect 332 11 334 13
rect 350 11 352 71
rect 366 11 368 71
rect 372 70 374 71
rect 372 68 376 70
rect 374 11 376 68
rect 390 11 392 71
rect 396 70 398 71
rect 396 68 400 70
rect 398 11 400 68
rect 414 11 416 71
rect 420 70 422 71
rect 420 68 424 70
rect 422 11 424 68
rect 438 11 440 71
rect 444 70 446 71
rect 444 68 448 70
rect 446 11 448 68
rect 463 11 465 71
rect 469 70 471 71
rect 469 68 473 70
rect 471 11 473 68
rect -172 4 -170 7
rect -164 4 -162 7
rect -140 4 -138 7
rect -117 4 -115 7
rect -94 4 -92 7
rect -86 4 -84 7
rect -70 4 -68 7
rect -62 4 -60 7
rect -6 4 -4 7
rect 2 4 4 7
rect 18 4 20 7
rect 34 4 36 7
rect 51 4 53 7
rect 57 4 59 7
rect 89 4 91 7
rect 113 4 115 7
rect 119 4 121 7
rect 137 4 139 7
rect 153 4 155 7
rect 161 4 163 7
rect 177 4 179 7
rect 185 4 187 7
rect 201 4 203 7
rect 209 4 211 7
rect 225 4 227 7
rect 233 4 235 7
rect 250 4 252 7
rect 258 4 260 7
rect 290 4 292 7
rect 296 4 298 7
rect 326 4 328 7
rect 332 4 334 7
rect 350 4 352 7
rect 366 4 368 7
rect 374 4 376 7
rect 390 4 392 7
rect 398 4 400 7
rect 414 4 416 7
rect 422 4 424 7
rect 438 4 440 7
rect 446 4 448 7
rect 463 4 465 7
rect 471 4 473 7
rect -180 -8 -178 -5
rect -158 -10 -156 -7
rect -132 -8 -130 -5
rect -126 -8 -124 -5
rect -118 -8 -116 -5
rect -88 -8 -86 -5
rect -80 -8 -78 -5
rect -74 -8 -72 -5
rect -56 -8 -54 -5
rect -180 -81 -178 -12
rect -32 -10 -30 -7
rect -10 -8 -8 -5
rect -4 -8 -2 -5
rect 4 -8 6 -5
rect 34 -8 36 -5
rect 42 -8 44 -5
rect 48 -8 50 -5
rect 82 -8 84 -5
rect 88 -8 90 -5
rect 96 -8 98 -5
rect 128 -8 130 -5
rect 136 -8 138 -5
rect 142 -8 144 -5
rect -158 -30 -156 -14
rect -158 -34 -155 -30
rect -158 -81 -156 -34
rect -132 -81 -130 -12
rect -126 -13 -124 -12
rect -127 -15 -124 -13
rect -127 -53 -125 -15
rect -118 -31 -116 -12
rect -118 -33 -114 -31
rect -127 -55 -122 -53
rect -124 -65 -122 -55
rect -124 -81 -122 -70
rect -116 -81 -114 -33
rect -88 -45 -86 -12
rect -80 -44 -78 -12
rect -90 -47 -86 -45
rect -82 -46 -78 -44
rect -90 -81 -88 -47
rect -82 -52 -80 -46
rect -82 -81 -80 -57
rect -74 -65 -72 -12
rect -74 -81 -72 -70
rect -56 -81 -54 -12
rect 164 -10 166 -7
rect 188 -8 190 -5
rect 206 -8 208 -5
rect 212 -8 214 -5
rect 220 -8 222 -5
rect 250 -8 252 -5
rect 258 -8 260 -5
rect 264 -8 266 -5
rect -32 -81 -30 -14
rect -10 -36 -8 -12
rect -4 -13 -2 -12
rect -9 -40 -8 -36
rect -10 -81 -8 -40
rect -5 -15 -2 -13
rect -5 -53 -3 -15
rect 4 -31 6 -12
rect 4 -33 8 -31
rect -5 -55 0 -53
rect -2 -65 0 -55
rect -2 -81 0 -70
rect 6 -81 8 -33
rect 34 -45 36 -12
rect 42 -44 44 -12
rect 32 -47 36 -45
rect 40 -46 44 -44
rect 32 -81 34 -47
rect 40 -52 42 -46
rect 40 -81 42 -57
rect 48 -65 50 -12
rect 82 -65 84 -12
rect 88 -44 90 -12
rect 88 -46 92 -44
rect 90 -52 92 -46
rect 96 -45 98 -12
rect 128 -31 130 -12
rect 136 -13 138 -12
rect 136 -15 139 -13
rect 126 -33 130 -31
rect 96 -47 100 -45
rect 48 -81 50 -70
rect 82 -81 84 -70
rect 90 -81 92 -57
rect 98 -81 100 -47
rect 126 -81 128 -33
rect 137 -53 139 -15
rect 134 -55 139 -53
rect 142 -36 144 -12
rect 290 -10 292 -7
rect 312 -8 314 -5
rect 349 -8 351 -5
rect 355 -8 357 -5
rect 363 -8 365 -5
rect 393 -8 395 -5
rect 401 -8 403 -5
rect 407 -8 409 -5
rect 142 -40 143 -36
rect 134 -65 136 -55
rect 134 -81 136 -70
rect 142 -81 144 -40
rect 164 -81 166 -14
rect 188 -81 190 -12
rect 206 -65 208 -12
rect 212 -44 214 -12
rect 212 -46 216 -44
rect 214 -52 216 -46
rect 220 -45 222 -12
rect 250 -31 252 -12
rect 258 -13 260 -12
rect 258 -15 261 -13
rect 248 -33 252 -31
rect 220 -47 224 -45
rect 206 -81 208 -70
rect 214 -81 216 -57
rect 222 -81 224 -47
rect 248 -81 250 -33
rect 259 -53 261 -15
rect 256 -55 261 -53
rect 256 -65 258 -55
rect 256 -81 258 -70
rect 264 -81 266 -12
rect 429 -10 431 -7
rect 453 -8 455 -5
rect 471 -8 473 -5
rect 477 -8 479 -5
rect 485 -8 487 -5
rect 515 -8 517 -5
rect 523 -8 525 -5
rect 529 -8 531 -5
rect 290 -21 292 -14
rect 289 -25 292 -21
rect 290 -81 292 -25
rect 312 -81 314 -12
rect 349 -65 351 -12
rect 355 -44 357 -12
rect 355 -46 359 -44
rect 357 -52 359 -46
rect 363 -45 365 -12
rect 393 -31 395 -12
rect 401 -13 403 -12
rect 401 -15 404 -13
rect 391 -33 395 -31
rect 363 -47 367 -45
rect 349 -81 351 -70
rect 357 -81 359 -57
rect 365 -81 367 -47
rect 391 -81 393 -33
rect 402 -53 404 -15
rect 399 -55 404 -53
rect 407 -36 409 -12
rect 558 -10 560 -7
rect 580 -8 582 -5
rect 407 -40 408 -36
rect 399 -65 401 -55
rect 399 -81 401 -70
rect 407 -81 409 -40
rect 429 -81 431 -14
rect 453 -81 455 -12
rect 471 -65 473 -12
rect 477 -44 479 -12
rect 477 -46 481 -44
rect 479 -52 481 -46
rect 485 -45 487 -12
rect 515 -31 517 -12
rect 523 -13 525 -12
rect 523 -15 526 -13
rect 513 -33 517 -31
rect 485 -47 489 -45
rect 471 -81 473 -70
rect 479 -81 481 -57
rect 487 -81 489 -47
rect 513 -81 515 -33
rect 524 -53 526 -15
rect 521 -55 526 -53
rect 521 -65 523 -55
rect 521 -81 523 -70
rect 529 -81 531 -12
rect 558 -30 560 -14
rect 557 -34 560 -30
rect 558 -81 560 -34
rect 580 -81 582 -12
rect -180 -92 -178 -89
rect -158 -92 -156 -89
rect -132 -92 -130 -89
rect -124 -92 -122 -89
rect -116 -92 -114 -89
rect -90 -92 -88 -89
rect -82 -92 -80 -89
rect -74 -92 -72 -89
rect -56 -92 -54 -89
rect -32 -92 -30 -89
rect -10 -92 -8 -89
rect -2 -92 0 -89
rect 6 -92 8 -89
rect 32 -92 34 -89
rect 40 -92 42 -89
rect 48 -92 50 -89
rect 82 -92 84 -89
rect 90 -92 92 -89
rect 98 -92 100 -89
rect 126 -92 128 -89
rect 134 -92 136 -89
rect 142 -92 144 -89
rect 164 -92 166 -89
rect 188 -92 190 -89
rect 206 -92 208 -89
rect 214 -92 216 -89
rect 222 -92 224 -89
rect 248 -92 250 -89
rect 256 -92 258 -89
rect 264 -92 266 -89
rect 290 -92 292 -89
rect 312 -92 314 -89
rect 349 -92 351 -89
rect 357 -92 359 -89
rect 365 -92 367 -89
rect 391 -92 393 -89
rect 399 -92 401 -89
rect 407 -92 409 -89
rect 429 -92 431 -89
rect 453 -92 455 -89
rect 471 -92 473 -89
rect 479 -92 481 -89
rect 487 -92 489 -89
rect 513 -92 515 -89
rect 521 -92 523 -89
rect 529 -92 531 -89
rect 558 -92 560 -89
rect 580 -92 582 -89
<< polycontact >>
rect -162 56 -158 60
rect -74 55 -70 59
rect 4 60 8 64
rect 14 41 18 45
rect 133 26 137 30
rect 149 14 153 18
rect 197 34 201 38
rect 221 20 225 24
rect 246 59 250 63
rect 346 26 350 30
rect 362 14 366 18
rect 410 14 414 18
rect 434 20 438 24
rect 459 59 463 63
rect -184 -54 -180 -50
rect -155 -34 -151 -30
rect -136 -34 -132 -30
rect -92 -29 -88 -25
rect -60 -70 -56 -66
rect -13 -40 -9 -36
rect 30 -29 34 -25
rect 98 -29 102 -25
rect 143 -40 147 -36
rect 222 -29 226 -25
rect 190 -70 194 -66
rect 266 -25 270 -21
rect 285 -25 289 -21
rect 314 -56 318 -52
rect 365 -29 369 -25
rect 408 -40 412 -36
rect 487 -29 491 -25
rect 455 -70 459 -66
rect 531 -34 535 -30
rect 553 -34 557 -30
rect 582 -56 586 -52
<< metal1 >>
rect -178 90 476 91
rect -178 89 13 90
rect -178 85 -176 89
rect -172 85 -168 89
rect -164 85 -160 89
rect -156 85 -145 89
rect -141 85 -137 89
rect -133 85 -122 89
rect -118 85 -114 89
rect -110 85 -100 89
rect -96 85 -92 89
rect -88 85 -84 89
rect -80 85 -74 89
rect -70 85 -66 89
rect -62 85 -58 89
rect -54 88 13 89
rect -54 85 -11 88
rect -178 84 -11 85
rect -7 84 3 88
rect 7 86 13 88
rect 17 86 21 90
rect 25 86 29 90
rect 33 86 37 90
rect 41 86 46 90
rect 50 86 54 90
rect 58 86 62 90
rect 66 86 84 90
rect 88 86 92 90
rect 96 86 108 90
rect 112 86 116 90
rect 120 86 124 90
rect 128 86 132 90
rect 136 86 140 90
rect 144 88 285 90
rect 144 86 148 88
rect 7 84 148 86
rect 152 84 162 88
rect 166 84 172 88
rect 176 84 186 88
rect 190 84 196 88
rect 200 84 210 88
rect 214 84 220 88
rect 224 84 234 88
rect 238 84 245 88
rect 249 84 259 88
rect 263 86 285 88
rect 289 86 293 90
rect 297 86 301 90
rect 305 86 321 90
rect 325 86 329 90
rect 333 86 337 90
rect 341 86 345 90
rect 349 86 353 90
rect 357 88 476 90
rect 357 86 361 88
rect 263 84 361 86
rect 365 84 375 88
rect 379 84 385 88
rect 389 84 399 88
rect 403 84 409 88
rect 413 84 423 88
rect 427 84 433 88
rect 437 84 447 88
rect 451 84 458 88
rect 462 84 472 88
rect -178 83 144 84
rect 148 83 357 84
rect 361 83 476 84
rect -161 79 -157 83
rect -137 79 -133 83
rect -122 79 -118 83
rect -99 79 -95 83
rect -59 79 -55 83
rect -175 49 -171 71
rect -145 60 -141 71
rect -158 56 -141 60
rect -175 45 -165 49
rect -169 11 -165 45
rect -145 11 -141 56
rect -114 44 -110 71
rect -85 59 -81 71
rect -11 79 -7 83
rect 13 79 17 83
rect 29 79 33 83
rect 46 79 50 83
rect 62 79 66 83
rect 84 79 88 83
rect 108 79 112 83
rect 124 79 128 83
rect 132 79 136 83
rect 148 79 152 83
rect 172 79 176 83
rect 196 79 200 83
rect 220 79 224 83
rect 245 79 249 83
rect 285 79 289 83
rect 301 79 305 83
rect 321 79 325 83
rect 337 79 341 83
rect 345 79 349 83
rect 361 79 365 83
rect 385 79 389 83
rect 409 79 413 83
rect 433 79 437 83
rect 458 79 462 83
rect -73 69 -69 71
rect -73 65 -63 69
rect -85 55 -74 59
rect -91 51 -81 55
rect -114 40 -106 44
rect -114 28 -110 40
rect -114 11 -110 23
rect -91 11 -87 51
rect -67 11 -63 65
rect -3 67 7 71
rect -3 45 1 67
rect -3 41 14 45
rect -3 11 1 41
rect 21 11 25 71
rect 37 65 41 71
rect 37 11 41 60
rect 54 38 58 71
rect 92 47 96 71
rect 92 42 97 47
rect 54 34 62 38
rect 54 15 58 34
rect 73 23 78 26
rect 54 11 64 15
rect 92 11 96 42
rect 116 30 120 71
rect 116 26 133 30
rect 116 15 120 26
rect 140 18 144 71
rect 156 67 166 71
rect 180 67 190 71
rect 204 67 214 71
rect 228 67 238 71
rect 253 67 263 71
rect 156 47 160 67
rect 156 43 164 47
rect 116 11 126 15
rect 140 14 149 18
rect 140 11 144 14
rect 156 11 160 43
rect 180 38 184 67
rect 180 34 197 38
rect 180 11 184 34
rect 204 24 208 67
rect 228 63 232 67
rect 228 59 246 63
rect 204 20 221 24
rect 204 11 208 20
rect 228 11 232 59
rect 253 39 257 67
rect 253 35 278 39
rect 253 11 257 35
rect 274 12 278 35
rect -177 3 -173 7
rect -161 3 -157 7
rect -137 3 -133 7
rect -122 3 -118 7
rect -99 3 -95 7
rect -83 3 -79 7
rect -75 3 -71 7
rect -59 3 -55 7
rect -11 3 -7 7
rect 5 3 9 7
rect 13 3 17 7
rect 29 3 33 7
rect 46 3 50 7
rect 84 3 88 7
rect 108 3 112 7
rect 132 3 136 7
rect 148 3 152 7
rect 164 3 168 7
rect 172 3 176 7
rect 188 3 192 7
rect 196 3 200 7
rect 212 3 216 7
rect 220 3 224 7
rect 236 3 240 7
rect 293 36 297 71
rect 293 32 301 36
rect 293 15 297 32
rect 329 30 333 71
rect 329 26 346 30
rect 329 15 333 26
rect 353 18 357 71
rect 369 67 379 71
rect 393 67 403 71
rect 417 67 427 71
rect 441 67 451 71
rect 466 67 476 71
rect 369 46 373 67
rect 369 42 377 46
rect 293 11 303 15
rect 329 11 339 15
rect 353 14 362 18
rect 353 11 357 14
rect 369 11 373 42
rect 393 18 397 67
rect 417 24 421 67
rect 441 63 445 67
rect 441 59 459 63
rect 417 20 434 24
rect 393 14 410 18
rect 393 11 397 14
rect 417 11 421 20
rect 441 11 445 59
rect 466 36 470 67
rect 466 32 489 36
rect 466 11 470 32
rect 245 3 249 7
rect 261 3 265 7
rect 285 3 289 7
rect 321 3 325 7
rect 345 3 349 7
rect 361 3 365 7
rect 377 3 381 7
rect 385 3 389 7
rect 401 3 405 7
rect 409 3 413 7
rect 425 3 429 7
rect 433 3 437 7
rect 449 3 453 7
rect 458 3 462 7
rect 474 3 478 7
rect -187 2 589 3
rect -187 -2 -185 2
rect -181 -2 -177 2
rect -49 -2 -37 2
rect -33 -2 -29 2
rect -25 -2 -15 2
rect 492 -2 510 2
rect 514 -2 518 2
rect 522 -2 532 2
rect 536 -2 553 2
rect 557 -2 561 2
rect 565 -2 575 2
rect 579 -2 583 2
rect 587 -2 589 2
rect -187 -4 589 -2
rect -185 -8 -181 -4
rect -155 -10 -151 -4
rect -196 -54 -184 -50
rect -177 -66 -173 -12
rect -137 -8 -133 -4
rect -115 -8 -111 -4
rect -93 -8 -89 -4
rect -71 -8 -67 -4
rect -61 -8 -57 -4
rect -29 -10 -25 -4
rect -163 -52 -159 -14
rect -123 -25 -119 -12
rect -123 -29 -92 -25
rect -151 -34 -146 -30
rect -140 -34 -136 -30
rect -162 -57 -159 -52
rect -177 -81 -173 -71
rect -163 -81 -159 -57
rect -137 -77 -117 -73
rect -137 -81 -133 -77
rect -121 -81 -117 -77
rect -113 -81 -109 -29
rect -85 -37 -81 -12
rect -90 -41 -81 -37
rect -95 -81 -91 -42
rect -71 -70 -60 -66
rect -87 -77 -67 -73
rect -87 -81 -83 -77
rect -71 -81 -67 -77
rect -53 -81 -49 -12
rect -15 -8 -11 -4
rect 7 -8 11 -4
rect 29 -8 33 -4
rect 51 -8 55 -4
rect 77 -8 81 -4
rect 99 -8 103 -4
rect 123 -8 127 -4
rect 145 -8 149 -4
rect 159 -10 163 -4
rect 191 -8 195 -4
rect -37 -52 -33 -14
rect -1 -25 3 -12
rect -1 -29 30 -25
rect -25 -40 -13 -36
rect -36 -57 -33 -52
rect -37 -81 -33 -57
rect -15 -77 5 -73
rect -15 -81 -11 -77
rect 1 -81 5 -77
rect 9 -81 13 -29
rect 37 -37 41 -12
rect 32 -41 41 -37
rect 91 -37 95 -12
rect 131 -25 135 -12
rect 102 -29 135 -25
rect 91 -41 100 -37
rect 27 -81 31 -42
rect 35 -77 55 -73
rect 35 -81 39 -77
rect 51 -81 55 -77
rect 77 -77 97 -73
rect 77 -81 81 -77
rect 93 -81 97 -77
rect 101 -81 105 -42
rect 121 -81 125 -29
rect 147 -40 159 -36
rect 167 -52 171 -14
rect 201 -8 205 -4
rect 223 -8 227 -4
rect 245 -8 249 -4
rect 267 -8 271 -4
rect 285 -10 289 -4
rect 315 -8 319 -4
rect 167 -57 170 -52
rect 129 -77 149 -73
rect 129 -81 133 -77
rect 145 -81 149 -77
rect 167 -81 171 -57
rect 183 -81 187 -12
rect 215 -37 219 -12
rect 253 -25 257 -12
rect 270 -25 273 -21
rect 279 -25 285 -21
rect 226 -29 257 -25
rect 215 -41 224 -37
rect 194 -70 205 -66
rect 201 -77 221 -73
rect 201 -81 205 -77
rect 217 -81 221 -77
rect 225 -81 229 -42
rect 243 -81 247 -29
rect 293 -52 297 -14
rect 344 -8 348 -4
rect 366 -8 370 -4
rect 388 -8 392 -4
rect 410 -8 414 -4
rect 424 -10 428 -4
rect 456 -8 460 -4
rect 293 -57 296 -52
rect 251 -77 271 -73
rect 251 -81 255 -77
rect 267 -81 271 -77
rect 293 -81 297 -57
rect 307 -66 311 -12
rect 358 -37 362 -12
rect 396 -25 400 -12
rect 369 -29 400 -25
rect 358 -41 367 -37
rect 318 -56 322 -52
rect 307 -81 311 -71
rect 344 -77 364 -73
rect 344 -81 348 -77
rect 360 -81 364 -77
rect 368 -81 372 -42
rect 386 -81 390 -29
rect 412 -40 424 -36
rect 432 -52 436 -14
rect 466 -8 470 -4
rect 488 -8 492 -4
rect 510 -8 514 -4
rect 532 -8 536 -4
rect 553 -10 557 -4
rect 583 -8 587 -4
rect 432 -57 435 -52
rect 394 -77 414 -73
rect 394 -81 398 -77
rect 410 -81 414 -77
rect 432 -81 436 -57
rect 448 -81 452 -12
rect 480 -37 484 -12
rect 518 -25 522 -12
rect 491 -29 522 -25
rect 480 -41 489 -37
rect 459 -70 470 -66
rect 466 -77 486 -73
rect 466 -81 470 -77
rect 482 -81 486 -77
rect 490 -81 494 -42
rect 508 -81 512 -29
rect 535 -34 541 -30
rect 547 -34 553 -30
rect 561 -52 565 -14
rect 561 -57 564 -52
rect 516 -77 536 -73
rect 516 -81 520 -77
rect 532 -81 536 -77
rect 561 -81 565 -57
rect 575 -66 579 -12
rect 586 -56 590 -52
rect 575 -81 579 -71
rect -185 -93 -181 -89
rect -155 -93 -151 -89
rect -129 -93 -125 -89
rect -79 -93 -75 -89
rect -61 -93 -57 -89
rect -29 -93 -25 -89
rect -7 -93 -3 -89
rect 43 -93 47 -89
rect 85 -93 89 -89
rect 137 -93 141 -89
rect 159 -93 163 -89
rect 191 -93 195 -89
rect 209 -93 213 -89
rect 259 -93 263 -89
rect 285 -93 289 -89
rect 315 -93 319 -89
rect 352 -93 356 -89
rect 402 -93 406 -89
rect 424 -93 428 -89
rect 456 -93 460 -89
rect 474 -93 478 -89
rect 524 -93 528 -89
rect 553 -93 557 -89
rect 583 -93 587 -89
rect -187 -95 589 -93
rect -187 -99 -185 -95
rect -181 -99 -177 -95
rect -173 -99 -163 -95
rect -159 -99 -155 -95
rect -151 -99 -137 -95
rect -133 -99 -129 -95
rect -125 -99 -121 -95
rect -117 -99 -113 -95
rect -109 -99 -95 -95
rect -91 -99 -87 -95
rect -83 -99 -79 -95
rect -75 -99 -71 -95
rect -67 -99 -37 -95
rect -33 -99 -29 -95
rect -25 -99 -15 -95
rect -11 -99 -7 -95
rect -3 -99 1 -95
rect 5 -99 9 -95
rect 13 -99 27 -95
rect 31 -99 35 -95
rect 39 -99 43 -95
rect 47 -99 51 -95
rect 55 -99 77 -95
rect 81 -99 85 -95
rect 89 -99 93 -95
rect 97 -99 101 -95
rect 105 -99 121 -95
rect 125 -99 129 -95
rect 133 -99 137 -95
rect 141 -99 145 -95
rect 149 -99 159 -95
rect 163 -99 167 -95
rect 171 -99 201 -95
rect 205 -99 209 -95
rect 213 -99 217 -95
rect 221 -99 225 -95
rect 229 -99 243 -95
rect 247 -99 251 -95
rect 255 -99 259 -95
rect 263 -99 267 -95
rect 271 -99 285 -95
rect 289 -99 293 -95
rect 297 -99 307 -95
rect 311 -99 315 -95
rect 319 -99 344 -95
rect 348 -99 352 -95
rect 356 -99 360 -95
rect 364 -99 368 -95
rect 372 -99 386 -95
rect 390 -99 394 -95
rect 398 -99 402 -95
rect 406 -99 410 -95
rect 414 -99 424 -95
rect 428 -99 432 -95
rect 436 -99 466 -95
rect 470 -99 474 -95
rect 478 -99 482 -95
rect 486 -99 490 -95
rect 494 -99 508 -95
rect 512 -99 516 -95
rect 520 -99 524 -95
rect 528 -99 532 -95
rect 536 -99 553 -95
rect 557 -99 561 -95
rect 565 -99 575 -95
rect 579 -99 583 -95
rect 587 -99 589 -95
rect -187 -101 589 -99
<< m2contact >>
rect -150 40 -145 45
rect -114 23 -109 28
rect 37 60 42 65
rect 25 52 30 57
rect 97 42 102 47
rect 62 34 67 39
rect 73 18 78 23
rect 164 42 169 47
rect 273 7 278 12
rect 301 32 306 37
rect 377 42 382 47
rect 489 32 494 37
rect -202 -55 -196 -50
rect -146 -34 -140 -29
rect -167 -57 -162 -52
rect -177 -71 -172 -66
rect -95 -42 -90 -37
rect -41 -57 -36 -52
rect -49 -71 -44 -66
rect 27 -42 32 -37
rect 100 -42 105 -37
rect 170 -57 175 -52
rect 178 -71 183 -66
rect 273 -25 279 -20
rect 224 -42 229 -37
rect 296 -57 301 -52
rect 367 -42 372 -37
rect 322 -56 328 -51
rect 306 -71 311 -66
rect 435 -57 440 -52
rect 443 -71 448 -66
rect 489 -42 494 -37
rect 541 -35 547 -30
rect 564 -57 569 -52
rect 590 -56 596 -51
rect 574 -71 579 -66
<< pm12contact >>
rect -177 23 -172 28
rect -122 48 -117 53
rect -99 48 -94 53
rect -138 14 -133 19
rect -84 40 -79 45
rect -12 59 -6 64
rect -60 38 -55 43
rect 4 26 9 31
rect 46 60 51 65
rect 29 29 34 34
rect 61 18 66 23
rect 84 18 89 23
rect 108 18 113 23
rect 123 18 128 23
rect 163 59 168 64
rect 172 16 177 21
rect 187 25 192 30
rect 211 34 216 39
rect 235 42 240 47
rect 285 60 290 65
rect 260 51 265 56
rect 300 42 305 47
rect 321 42 326 47
rect 336 18 341 23
rect 376 59 381 64
rect 385 18 390 23
rect 400 21 405 26
rect 424 32 429 37
rect 448 42 453 47
rect 473 51 478 56
rect -121 -42 -116 -37
rect -126 -70 -121 -65
rect -84 -57 -79 -52
rect -76 -70 -71 -65
rect -30 -41 -25 -36
rect 1 -42 6 -37
rect -4 -70 1 -65
rect 38 -57 43 -52
rect 89 -57 94 -52
rect 46 -70 51 -65
rect 81 -70 86 -65
rect 128 -42 133 -37
rect 159 -41 164 -36
rect 133 -70 138 -65
rect 213 -57 218 -52
rect 205 -70 210 -65
rect 250 -42 255 -37
rect 255 -70 260 -65
rect 356 -57 361 -52
rect 348 -70 353 -65
rect 393 -42 398 -37
rect 424 -41 429 -36
rect 398 -70 403 -65
rect 478 -57 483 -52
rect 470 -70 475 -65
rect 515 -42 520 -37
rect 520 -70 525 -65
<< metal2 >>
rect -133 53 -128 56
rect 42 60 46 64
rect 51 60 163 64
rect 168 60 285 64
rect 290 60 376 64
rect -133 48 -122 53
rect -117 48 -99 52
rect -145 40 -84 44
rect -12 43 -7 59
rect 30 51 260 55
rect 265 51 473 55
rect -55 38 -7 43
rect 95 42 97 47
rect 102 42 105 47
rect 110 42 112 47
rect 169 43 235 47
rect 305 42 310 47
rect 317 42 321 47
rect 382 43 448 47
rect -172 23 -114 27
rect -133 14 -29 18
rect -12 -11 -7 38
rect 67 34 211 38
rect 9 26 21 30
rect -145 -16 -7 -11
rect -145 -29 -140 -16
rect -116 -41 -95 -37
rect -90 -41 -30 -37
rect 17 -37 21 26
rect 306 33 424 37
rect 29 21 33 29
rect 192 25 194 30
rect 199 25 200 30
rect 66 18 73 22
rect 78 18 84 22
rect 89 18 108 22
rect 128 18 172 22
rect 177 17 336 21
rect 341 18 385 22
rect 405 21 408 26
rect 489 27 494 32
rect 489 23 546 27
rect 29 10 33 16
rect 29 6 116 10
rect 112 -37 116 6
rect 273 -20 278 7
rect 379 -14 383 18
rect 6 -41 27 -37
rect 105 -41 128 -37
rect 379 -37 383 -19
rect 542 -30 546 23
rect 164 -41 224 -37
rect 229 -41 250 -37
rect -202 -50 -196 -44
rect 372 -41 393 -37
rect 429 -41 489 -37
rect 494 -41 515 -37
rect 322 -51 328 -44
rect -162 -56 -84 -52
rect -36 -56 38 -52
rect 94 -56 170 -52
rect 218 -56 296 -52
rect 590 -51 596 -44
rect 361 -56 435 -52
rect 483 -56 564 -52
rect -172 -70 -126 -66
rect -121 -70 -76 -66
rect -44 -70 -4 -66
rect 1 -70 46 -66
rect 86 -70 133 -66
rect 138 -70 178 -66
rect 210 -70 255 -66
rect 260 -70 306 -66
rect 353 -70 398 -66
rect 403 -70 443 -66
rect 475 -70 520 -66
rect 525 -70 574 -66
<< m3contact >>
rect -135 56 -128 62
rect 105 42 110 47
rect 310 42 317 47
rect -29 14 -22 21
rect -202 -44 -196 -38
rect 194 25 199 30
rect 408 21 413 29
rect 378 -19 384 -14
rect 322 -44 328 -38
rect 590 -44 596 -38
<< m123contact >>
rect 28 16 33 21
<< metal3 >>
rect -128 56 -37 61
rect -42 -14 -37 56
rect 110 42 310 47
rect 199 29 413 30
rect 199 25 408 29
rect -22 16 28 21
rect -42 -19 378 -14
rect -196 -44 322 -38
rect 328 -44 590 -38
<< labels >>
rlabel polycontact 4 60 8 64 1 RST
rlabel metal1 10 83 10 91 1 VDD
rlabel metal1 10 -5 10 3 1 GND
rlabel pm12contact 187 25 192 30 1 REQ
rlabel metal1 73 23 78 26 1 T
rlabel pm12contact -136 16 -136 16 1 s1
rlabel metal1 -175 57 -171 59 1 RED
rlabel metal1 -145 56 -141 60 1 GREEN
rlabel metal1 -91 48 -87 51 1 YELLOW
rlabel metal1 -67 37 -63 41 1 S
<< end >>
